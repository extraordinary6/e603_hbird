 /*                                                                      
  *  Copyright (c) 2018-2025 Nuclei System Technology, Inc.       
  *  All rights reserved.                                                
  */                                                                     
`include "global.v"
module e603_sram_icb_ctrl #(
    parameter ECC = 0,
    parameter CS_W = 1,
    parameter DW = 32,
    parameter MW = 4,
    parameter AW = 32,
    parameter AW_LSB = 3,
    parameter RAM_DW = DW,
    parameter RAM_MW = MW,
    parameter DELAY_WIDTH=9,
    parameter USR_W = 3 
)(
  input  [DELAY_WIDTH-1:0] delay_select,
  output sram_ctrl_active,
  input  tcm_cgstop,
  input  stall_uop_cmd,
  input  i_icb_cmd_valid, 
  output i_icb_cmd_ready, 
  input  i_icb_cmd_read,  
  input  [AW-1:0] i_icb_cmd_addr, 
  input  [DW-1:0] i_icb_cmd_wdata, 
  input  [MW-1:0] i_icb_cmd_wmask, 
  input  [USR_W-1:0] i_icb_cmd_usr, 
  output i_icb_rsp_valid, 
  input  i_icb_rsp_ready, 
  output [DW-1:0] i_icb_rsp_rdata, 
  output [USR_W-1:0] i_icb_rsp_usr, 
  output i_icb_rsp_err, 
  output [CS_W-1:0]      ram_cs,  
  output [AW-AW_LSB-1:0] ram_addr, 
  output [CS_W-1:0]      ram_we,  
  output [RAM_MW-1:0] ram_wem,
  output [RAM_DW-1:0] ram_din,          
  input  [RAM_DW-1:0] ram_dout,
  output          clk_ram,
  input  clkgate_bypass,
  input  clk,
  input  rst_n
  );
  wire  byp_icb_cmd_valid;
  wire  byp_icb_cmd_ready;
  wire  byp_icb_cmd_read;
  wire  [AW-1:0] byp_icb_cmd_addr; 
  wire  [DW-1:0] byp_icb_cmd_wdata; 
  wire  [MW-1:0] byp_icb_cmd_wmask; 
  wire  [USR_W-1:0] byp_icb_cmd_usr; 
e603_ddr_icb_cmd_delay #(
    .DW (DW),
    .MW (MW),
    .AW (AW),
    .USR_W (USR_W) 
)u_icb_cmd_delay(
  .i_icb_cmd_valid      (i_icb_cmd_valid ), 
  .i_icb_cmd_ready      (i_icb_cmd_ready ), 
  .i_icb_cmd_read       (i_icb_cmd_read  ),  
  .i_icb_cmd_addr       (i_icb_cmd_addr  ), 
  .i_icb_cmd_wdata      (i_icb_cmd_wdata ), 
  .i_icb_cmd_wmask      (i_icb_cmd_wmask ), 
  .i_icb_cmd_usr        (i_icb_cmd_usr   ), 
  .o_icb_cmd_valid      (byp_icb_cmd_valid ), 
  .o_icb_cmd_ready      (byp_icb_cmd_ready ), 
  .o_icb_cmd_read       (byp_icb_cmd_read  ),  
  .o_icb_cmd_addr       (byp_icb_cmd_addr  ), 
  .o_icb_cmd_wdata      (byp_icb_cmd_wdata ), 
  .o_icb_cmd_wmask      (byp_icb_cmd_wmask ), 
  .o_icb_cmd_usr        (byp_icb_cmd_usr   ), 
  .delay_select         (delay_select),
  .clkgate_bypass       (clkgate_bypass  ),
  .clk                  (clk             ),
  .rst_n                (rst_n           )
  );
  wire sram_active;
generate
if (ECC == 0)
begin: noecc
  e603_1cyc_sram_ctrl #(
      .CS_W   (CS_W),
      .DW     (DW),
      .AW     (AW),
      .MW     (MW),
      .AW_LSB (AW_LSB),
      .USR_W  (USR_W) 
  ) u_1cyc_sram_ctrl(
     .sram_ctrl_active (sram_active),
     .tcm_cgstop       (tcm_cgstop),
     .stall_uop_cmd (stall_uop_cmd),
     .uop_cmd_valid (byp_icb_cmd_valid),
     .uop_cmd_ready (byp_icb_cmd_ready),
     .uop_cmd_read  (byp_icb_cmd_read ),
     .uop_cmd_addr  (byp_icb_cmd_addr ), 
     .uop_cmd_size  (2'b0             ), 
     .uop_cmd_wdata (byp_icb_cmd_wdata), 
     .uop_cmd_wmask (byp_icb_cmd_wmask), 
     .uop_cmd_usr   (byp_icb_cmd_usr  ),
     .uop_rsp_valid (i_icb_rsp_valid),
     .uop_rsp_ready (i_icb_rsp_ready),
     .uop_rsp_err   (               ),
     .uop_rsp_rdata (i_icb_rsp_rdata),
     .uop_rsp_usr   (i_icb_rsp_usr  ),
     .ram_cs   (ram_cs  ),  
     .ram_addr (ram_addr), 
     .ram_wem  (ram_wem ),
     .ram_we   (ram_we  ),
     .ram_din  (ram_din ),          
     .ram_dout (ram_dout),
     .clk_ram  (clk_ram ),
     .clkgate_bypass(clkgate_bypass  ),
     .clk  (clk  ),
     .rst_n(rst_n)  
    );
  assign i_icb_rsp_err = 1'b0;
end else begin : ecc
  e603_ilm_icb2sram_ecc u_ecc_icb_ctrl(
     .sram_wq_active (),
     .sram_ctrl_active (sram_active),
     .csr_ena_ecc_prot (1'b0),
     .csr_ena_ecc_chck (1'b0),
     .csr_ena_ecc_excp (1'b0),
     .csr_ecc_code_en  (1'b0),
     .csr_ecc_code     (8'b0),
     .ecc_dberr_pulse    (),
     .ecc_sberr_pulse    (),
     .stall_uop_cmd   (stall_uop_cmd),
     .icb_cmd_valid (byp_icb_cmd_valid),
     .icb_cmd_ready (byp_icb_cmd_ready),
     .icb_cmd_read  (byp_icb_cmd_read ),
     .icb_cmd_addr  (byp_icb_cmd_addr ), 
     .icb_cmd_wdata (byp_icb_cmd_wdata), 
     .icb_cmd_wmask (byp_icb_cmd_wmask), 
     .icb_cmd_size  (2'b11 ), 
     .icb_cmd_dmode (1'b0 ), 
     .icb_rsp_valid (i_icb_rsp_valid),
     .icb_rsp_ready (i_icb_rsp_ready),
     .icb_rsp_rdata (i_icb_rsp_rdata),
     .icb_rsp_err   (i_icb_rsp_err  ),
     .icb_rsp_eccerr(               ),
     .ram_dmode   (),  
     .ram_cs   (ram_cs  ),  
     .ram_addr (ram_addr), 
     .ram_we   (ram_we  ),
     .ram_wem  (ram_wem ),
     .ram_din  (ram_din ),          
     .ram_dout (ram_dout),
     .ram_clk  (clk_ram ),
     .clkgate_bypass       (clkgate_bypass),
     .clk  (clk  ),
     .rst_n(rst_n)  
    );
  assign i_icb_rsp_usr = {USR_W{1'b0}};
end
endgenerate
  assign sram_ctrl_active = 
                       i_icb_cmd_valid 
                     | byp_icb_cmd_valid 
                     | sram_active  
                     | i_icb_rsp_valid 
                     ;
endmodule
module e603_ddr_icb_cmd_delay #(
    parameter DW = 32,
    parameter MW = 4,
    parameter AW = 32,
    parameter USR_W = 3 
)(
  input  i_icb_cmd_valid, 
  output i_icb_cmd_ready, 
  input  i_icb_cmd_read,  
  input  [AW-1:0] i_icb_cmd_addr, 
  input  [DW-1:0] i_icb_cmd_wdata, 
  input  [MW-1:0] i_icb_cmd_wmask, 
  input  [USR_W-1:0] i_icb_cmd_usr, 
  output o_icb_cmd_valid, 
  input  o_icb_cmd_ready, 
  output o_icb_cmd_read,  
  output [AW-1:0] o_icb_cmd_addr, 
  output [DW-1:0] o_icb_cmd_wdata, 
  output [MW-1:0] o_icb_cmd_wmask, 
  output [USR_W-1:0] o_icb_cmd_usr, 
  input [9-1:0] delay_select,
  input  clkgate_bypass,
  input  clk,
  input  rst_n
  );
  wire  byp_icb_cmd_valid;
  wire  byp_icb_cmd_ready;
  wire  byp_icb_cmd_read;
  wire  [AW-1:0] byp_icb_cmd_addr; 
  wire  [DW-1:0] byp_icb_cmd_wdata; 
  wire  [MW-1:0] byp_icb_cmd_wmask; 
  wire  [USR_W-1:0] byp_icb_cmd_usr; 
  localparam BUF_CMD_PACK_W = (AW+DW+MW+USR_W+1);
  wire [BUF_CMD_PACK_W-1:0] byp_icb_cmd_o_pack;
  wire [BUF_CMD_PACK_W-1:0] byp_icb_cmd_i_pack =  {
                      i_icb_cmd_read, 
                      i_icb_cmd_addr, 
                      i_icb_cmd_wdata, 
                      i_icb_cmd_wmask, 
                      i_icb_cmd_usr  
                    };
  assign {
                      byp_icb_cmd_read, 
                      byp_icb_cmd_addr, 
                      byp_icb_cmd_wdata, 
                      byp_icb_cmd_wmask, 
                      byp_icb_cmd_usr  
                    } = byp_icb_cmd_o_pack;
`ifdef SYNTHESIS 
  e603_gnrl_bypbuf # (
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_byp_icb_cmd_buf(
    .i_vld(i_icb_cmd_valid), 
    .i_rdy(i_icb_cmd_ready), 
    .i_dat(byp_icb_cmd_i_pack),
    .o_vld(byp_icb_cmd_valid), 
    .o_rdy(byp_icb_cmd_ready), 
    .o_dat(byp_icb_cmd_o_pack),
    .fifo_o_vld(),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
`else 
`ifdef NO_CCT_DDR_LATENCY
  e603_gnrl_bypbuf # (
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_byp_icb_cmd_buf(
    .i_vld(i_icb_cmd_valid), 
    .i_rdy(i_icb_cmd_ready), 
    .i_dat(byp_icb_cmd_i_pack),
    .o_vld(byp_icb_cmd_valid), 
    .o_rdy(byp_icb_cmd_ready), 
    .o_dat(byp_icb_cmd_o_pack),
    .fifo_o_vld(),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
`else
  wire [511:0] delay_stage_select = 512'b1 << delay_select;
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_0;
  wire     tmp_icb_cmd_valid_0;
  wire     tmp_icb_cmd_ready_0;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_0 (
    .i_vld(i_icb_cmd_valid), 
    .i_rdy(i_icb_cmd_ready), 
    .i_dat(byp_icb_cmd_i_pack),
    .o_vld(tmp_icb_cmd_valid_0), 
    .o_rdy(delay_stage_select[0] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_0), 
    .o_dat(tmp_icb_cmd_pack_0),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_1;
  wire     tmp_icb_cmd_valid_1;
  wire     tmp_icb_cmd_ready_1;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_1 (
    .i_vld(tmp_icb_cmd_valid_0), 
    .i_rdy(tmp_icb_cmd_ready_0), 
    .i_dat(tmp_icb_cmd_pack_0),
    .o_vld(tmp_icb_cmd_valid_1), 
    .o_rdy(delay_stage_select[1] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_1), 
    .o_dat(tmp_icb_cmd_pack_1),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_2;
  wire     tmp_icb_cmd_valid_2;
  wire     tmp_icb_cmd_ready_2;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_2 (
    .i_vld(tmp_icb_cmd_valid_1), 
    .i_rdy(tmp_icb_cmd_ready_1), 
    .i_dat(tmp_icb_cmd_pack_1),
    .o_vld(tmp_icb_cmd_valid_2), 
    .o_rdy(delay_stage_select[2] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_2), 
    .o_dat(tmp_icb_cmd_pack_2),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_3;
  wire     tmp_icb_cmd_valid_3;
  wire     tmp_icb_cmd_ready_3;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_3 (
    .i_vld(tmp_icb_cmd_valid_2), 
    .i_rdy(tmp_icb_cmd_ready_2), 
    .i_dat(tmp_icb_cmd_pack_2),
    .o_vld(tmp_icb_cmd_valid_3), 
    .o_rdy(delay_stage_select[3] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_3), 
    .o_dat(tmp_icb_cmd_pack_3),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_4;
  wire     tmp_icb_cmd_valid_4;
  wire     tmp_icb_cmd_ready_4;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_4 (
    .i_vld(tmp_icb_cmd_valid_3), 
    .i_rdy(tmp_icb_cmd_ready_3), 
    .i_dat(tmp_icb_cmd_pack_3),
    .o_vld(tmp_icb_cmd_valid_4), 
    .o_rdy(delay_stage_select[4] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_4), 
    .o_dat(tmp_icb_cmd_pack_4),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_5;
  wire     tmp_icb_cmd_valid_5;
  wire     tmp_icb_cmd_ready_5;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_5 (
    .i_vld(tmp_icb_cmd_valid_4), 
    .i_rdy(tmp_icb_cmd_ready_4), 
    .i_dat(tmp_icb_cmd_pack_4),
    .o_vld(tmp_icb_cmd_valid_5), 
    .o_rdy(delay_stage_select[5] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_5), 
    .o_dat(tmp_icb_cmd_pack_5),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_6;
  wire     tmp_icb_cmd_valid_6;
  wire     tmp_icb_cmd_ready_6;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_6 (
    .i_vld(tmp_icb_cmd_valid_5), 
    .i_rdy(tmp_icb_cmd_ready_5), 
    .i_dat(tmp_icb_cmd_pack_5),
    .o_vld(tmp_icb_cmd_valid_6), 
    .o_rdy(delay_stage_select[6] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_6), 
    .o_dat(tmp_icb_cmd_pack_6),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_7;
  wire     tmp_icb_cmd_valid_7;
  wire     tmp_icb_cmd_ready_7;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_7 (
    .i_vld(tmp_icb_cmd_valid_6), 
    .i_rdy(tmp_icb_cmd_ready_6), 
    .i_dat(tmp_icb_cmd_pack_6),
    .o_vld(tmp_icb_cmd_valid_7), 
    .o_rdy(delay_stage_select[7] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_7), 
    .o_dat(tmp_icb_cmd_pack_7),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_8;
  wire     tmp_icb_cmd_valid_8;
  wire     tmp_icb_cmd_ready_8;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_8 (
    .i_vld(tmp_icb_cmd_valid_7), 
    .i_rdy(tmp_icb_cmd_ready_7), 
    .i_dat(tmp_icb_cmd_pack_7),
    .o_vld(tmp_icb_cmd_valid_8), 
    .o_rdy(delay_stage_select[8] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_8), 
    .o_dat(tmp_icb_cmd_pack_8),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_9;
  wire     tmp_icb_cmd_valid_9;
  wire     tmp_icb_cmd_ready_9;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_9 (
    .i_vld(tmp_icb_cmd_valid_8), 
    .i_rdy(tmp_icb_cmd_ready_8), 
    .i_dat(tmp_icb_cmd_pack_8),
    .o_vld(tmp_icb_cmd_valid_9), 
    .o_rdy(delay_stage_select[9] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_9), 
    .o_dat(tmp_icb_cmd_pack_9),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_10;
  wire     tmp_icb_cmd_valid_10;
  wire     tmp_icb_cmd_ready_10;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_10 (
    .i_vld(tmp_icb_cmd_valid_9), 
    .i_rdy(tmp_icb_cmd_ready_9), 
    .i_dat(tmp_icb_cmd_pack_9),
    .o_vld(tmp_icb_cmd_valid_10), 
    .o_rdy(delay_stage_select[10] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_10), 
    .o_dat(tmp_icb_cmd_pack_10),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_11;
  wire     tmp_icb_cmd_valid_11;
  wire     tmp_icb_cmd_ready_11;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_11 (
    .i_vld(tmp_icb_cmd_valid_10), 
    .i_rdy(tmp_icb_cmd_ready_10), 
    .i_dat(tmp_icb_cmd_pack_10),
    .o_vld(tmp_icb_cmd_valid_11), 
    .o_rdy(delay_stage_select[11] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_11), 
    .o_dat(tmp_icb_cmd_pack_11),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_12;
  wire     tmp_icb_cmd_valid_12;
  wire     tmp_icb_cmd_ready_12;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_12 (
    .i_vld(tmp_icb_cmd_valid_11), 
    .i_rdy(tmp_icb_cmd_ready_11), 
    .i_dat(tmp_icb_cmd_pack_11),
    .o_vld(tmp_icb_cmd_valid_12), 
    .o_rdy(delay_stage_select[12] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_12), 
    .o_dat(tmp_icb_cmd_pack_12),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_13;
  wire     tmp_icb_cmd_valid_13;
  wire     tmp_icb_cmd_ready_13;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_13 (
    .i_vld(tmp_icb_cmd_valid_12), 
    .i_rdy(tmp_icb_cmd_ready_12), 
    .i_dat(tmp_icb_cmd_pack_12),
    .o_vld(tmp_icb_cmd_valid_13), 
    .o_rdy(delay_stage_select[13] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_13), 
    .o_dat(tmp_icb_cmd_pack_13),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_14;
  wire     tmp_icb_cmd_valid_14;
  wire     tmp_icb_cmd_ready_14;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_14 (
    .i_vld(tmp_icb_cmd_valid_13), 
    .i_rdy(tmp_icb_cmd_ready_13), 
    .i_dat(tmp_icb_cmd_pack_13),
    .o_vld(tmp_icb_cmd_valid_14), 
    .o_rdy(delay_stage_select[14] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_14), 
    .o_dat(tmp_icb_cmd_pack_14),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_15;
  wire     tmp_icb_cmd_valid_15;
  wire     tmp_icb_cmd_ready_15;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_15 (
    .i_vld(tmp_icb_cmd_valid_14), 
    .i_rdy(tmp_icb_cmd_ready_14), 
    .i_dat(tmp_icb_cmd_pack_14),
    .o_vld(tmp_icb_cmd_valid_15), 
    .o_rdy(delay_stage_select[15] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_15), 
    .o_dat(tmp_icb_cmd_pack_15),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_16;
  wire     tmp_icb_cmd_valid_16;
  wire     tmp_icb_cmd_ready_16;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_16 (
    .i_vld(tmp_icb_cmd_valid_15), 
    .i_rdy(tmp_icb_cmd_ready_15), 
    .i_dat(tmp_icb_cmd_pack_15),
    .o_vld(tmp_icb_cmd_valid_16), 
    .o_rdy(delay_stage_select[16] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_16), 
    .o_dat(tmp_icb_cmd_pack_16),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_17;
  wire     tmp_icb_cmd_valid_17;
  wire     tmp_icb_cmd_ready_17;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_17 (
    .i_vld(tmp_icb_cmd_valid_16), 
    .i_rdy(tmp_icb_cmd_ready_16), 
    .i_dat(tmp_icb_cmd_pack_16),
    .o_vld(tmp_icb_cmd_valid_17), 
    .o_rdy(delay_stage_select[17] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_17), 
    .o_dat(tmp_icb_cmd_pack_17),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_18;
  wire     tmp_icb_cmd_valid_18;
  wire     tmp_icb_cmd_ready_18;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_18 (
    .i_vld(tmp_icb_cmd_valid_17), 
    .i_rdy(tmp_icb_cmd_ready_17), 
    .i_dat(tmp_icb_cmd_pack_17),
    .o_vld(tmp_icb_cmd_valid_18), 
    .o_rdy(delay_stage_select[18] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_18), 
    .o_dat(tmp_icb_cmd_pack_18),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_19;
  wire     tmp_icb_cmd_valid_19;
  wire     tmp_icb_cmd_ready_19;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_19 (
    .i_vld(tmp_icb_cmd_valid_18), 
    .i_rdy(tmp_icb_cmd_ready_18), 
    .i_dat(tmp_icb_cmd_pack_18),
    .o_vld(tmp_icb_cmd_valid_19), 
    .o_rdy(delay_stage_select[19] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_19), 
    .o_dat(tmp_icb_cmd_pack_19),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_20;
  wire     tmp_icb_cmd_valid_20;
  wire     tmp_icb_cmd_ready_20;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_20 (
    .i_vld(tmp_icb_cmd_valid_19), 
    .i_rdy(tmp_icb_cmd_ready_19), 
    .i_dat(tmp_icb_cmd_pack_19),
    .o_vld(tmp_icb_cmd_valid_20), 
    .o_rdy(delay_stage_select[20] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_20), 
    .o_dat(tmp_icb_cmd_pack_20),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_21;
  wire     tmp_icb_cmd_valid_21;
  wire     tmp_icb_cmd_ready_21;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_21 (
    .i_vld(tmp_icb_cmd_valid_20), 
    .i_rdy(tmp_icb_cmd_ready_20), 
    .i_dat(tmp_icb_cmd_pack_20),
    .o_vld(tmp_icb_cmd_valid_21), 
    .o_rdy(delay_stage_select[21] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_21), 
    .o_dat(tmp_icb_cmd_pack_21),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_22;
  wire     tmp_icb_cmd_valid_22;
  wire     tmp_icb_cmd_ready_22;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_22 (
    .i_vld(tmp_icb_cmd_valid_21), 
    .i_rdy(tmp_icb_cmd_ready_21), 
    .i_dat(tmp_icb_cmd_pack_21),
    .o_vld(tmp_icb_cmd_valid_22), 
    .o_rdy(delay_stage_select[22] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_22), 
    .o_dat(tmp_icb_cmd_pack_22),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_23;
  wire     tmp_icb_cmd_valid_23;
  wire     tmp_icb_cmd_ready_23;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_23 (
    .i_vld(tmp_icb_cmd_valid_22), 
    .i_rdy(tmp_icb_cmd_ready_22), 
    .i_dat(tmp_icb_cmd_pack_22),
    .o_vld(tmp_icb_cmd_valid_23), 
    .o_rdy(delay_stage_select[23] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_23), 
    .o_dat(tmp_icb_cmd_pack_23),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_24;
  wire     tmp_icb_cmd_valid_24;
  wire     tmp_icb_cmd_ready_24;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_24 (
    .i_vld(tmp_icb_cmd_valid_23), 
    .i_rdy(tmp_icb_cmd_ready_23), 
    .i_dat(tmp_icb_cmd_pack_23),
    .o_vld(tmp_icb_cmd_valid_24), 
    .o_rdy(delay_stage_select[24] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_24), 
    .o_dat(tmp_icb_cmd_pack_24),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_25;
  wire     tmp_icb_cmd_valid_25;
  wire     tmp_icb_cmd_ready_25;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_25 (
    .i_vld(tmp_icb_cmd_valid_24), 
    .i_rdy(tmp_icb_cmd_ready_24), 
    .i_dat(tmp_icb_cmd_pack_24),
    .o_vld(tmp_icb_cmd_valid_25), 
    .o_rdy(delay_stage_select[25] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_25), 
    .o_dat(tmp_icb_cmd_pack_25),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_26;
  wire     tmp_icb_cmd_valid_26;
  wire     tmp_icb_cmd_ready_26;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_26 (
    .i_vld(tmp_icb_cmd_valid_25), 
    .i_rdy(tmp_icb_cmd_ready_25), 
    .i_dat(tmp_icb_cmd_pack_25),
    .o_vld(tmp_icb_cmd_valid_26), 
    .o_rdy(delay_stage_select[26] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_26), 
    .o_dat(tmp_icb_cmd_pack_26),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_27;
  wire     tmp_icb_cmd_valid_27;
  wire     tmp_icb_cmd_ready_27;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_27 (
    .i_vld(tmp_icb_cmd_valid_26), 
    .i_rdy(tmp_icb_cmd_ready_26), 
    .i_dat(tmp_icb_cmd_pack_26),
    .o_vld(tmp_icb_cmd_valid_27), 
    .o_rdy(delay_stage_select[27] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_27), 
    .o_dat(tmp_icb_cmd_pack_27),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_28;
  wire     tmp_icb_cmd_valid_28;
  wire     tmp_icb_cmd_ready_28;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_28 (
    .i_vld(tmp_icb_cmd_valid_27), 
    .i_rdy(tmp_icb_cmd_ready_27), 
    .i_dat(tmp_icb_cmd_pack_27),
    .o_vld(tmp_icb_cmd_valid_28), 
    .o_rdy(delay_stage_select[28] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_28), 
    .o_dat(tmp_icb_cmd_pack_28),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_29;
  wire     tmp_icb_cmd_valid_29;
  wire     tmp_icb_cmd_ready_29;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_29 (
    .i_vld(tmp_icb_cmd_valid_28), 
    .i_rdy(tmp_icb_cmd_ready_28), 
    .i_dat(tmp_icb_cmd_pack_28),
    .o_vld(tmp_icb_cmd_valid_29), 
    .o_rdy(delay_stage_select[29] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_29), 
    .o_dat(tmp_icb_cmd_pack_29),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_30;
  wire     tmp_icb_cmd_valid_30;
  wire     tmp_icb_cmd_ready_30;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_30 (
    .i_vld(tmp_icb_cmd_valid_29), 
    .i_rdy(tmp_icb_cmd_ready_29), 
    .i_dat(tmp_icb_cmd_pack_29),
    .o_vld(tmp_icb_cmd_valid_30), 
    .o_rdy(delay_stage_select[30] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_30), 
    .o_dat(tmp_icb_cmd_pack_30),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_31;
  wire     tmp_icb_cmd_valid_31;
  wire     tmp_icb_cmd_ready_31;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_31 (
    .i_vld(tmp_icb_cmd_valid_30), 
    .i_rdy(tmp_icb_cmd_ready_30), 
    .i_dat(tmp_icb_cmd_pack_30),
    .o_vld(tmp_icb_cmd_valid_31), 
    .o_rdy(delay_stage_select[31] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_31), 
    .o_dat(tmp_icb_cmd_pack_31),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_32;
  wire     tmp_icb_cmd_valid_32;
  wire     tmp_icb_cmd_ready_32;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_32 (
    .i_vld(tmp_icb_cmd_valid_31), 
    .i_rdy(tmp_icb_cmd_ready_31), 
    .i_dat(tmp_icb_cmd_pack_31),
    .o_vld(tmp_icb_cmd_valid_32), 
    .o_rdy(delay_stage_select[32] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_32), 
    .o_dat(tmp_icb_cmd_pack_32),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_33;
  wire     tmp_icb_cmd_valid_33;
  wire     tmp_icb_cmd_ready_33;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_33 (
    .i_vld(tmp_icb_cmd_valid_32), 
    .i_rdy(tmp_icb_cmd_ready_32), 
    .i_dat(tmp_icb_cmd_pack_32),
    .o_vld(tmp_icb_cmd_valid_33), 
    .o_rdy(delay_stage_select[33] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_33), 
    .o_dat(tmp_icb_cmd_pack_33),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_34;
  wire     tmp_icb_cmd_valid_34;
  wire     tmp_icb_cmd_ready_34;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_34 (
    .i_vld(tmp_icb_cmd_valid_33), 
    .i_rdy(tmp_icb_cmd_ready_33), 
    .i_dat(tmp_icb_cmd_pack_33),
    .o_vld(tmp_icb_cmd_valid_34), 
    .o_rdy(delay_stage_select[34] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_34), 
    .o_dat(tmp_icb_cmd_pack_34),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_35;
  wire     tmp_icb_cmd_valid_35;
  wire     tmp_icb_cmd_ready_35;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_35 (
    .i_vld(tmp_icb_cmd_valid_34), 
    .i_rdy(tmp_icb_cmd_ready_34), 
    .i_dat(tmp_icb_cmd_pack_34),
    .o_vld(tmp_icb_cmd_valid_35), 
    .o_rdy(delay_stage_select[35] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_35), 
    .o_dat(tmp_icb_cmd_pack_35),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_36;
  wire     tmp_icb_cmd_valid_36;
  wire     tmp_icb_cmd_ready_36;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_36 (
    .i_vld(tmp_icb_cmd_valid_35), 
    .i_rdy(tmp_icb_cmd_ready_35), 
    .i_dat(tmp_icb_cmd_pack_35),
    .o_vld(tmp_icb_cmd_valid_36), 
    .o_rdy(delay_stage_select[36] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_36), 
    .o_dat(tmp_icb_cmd_pack_36),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_37;
  wire     tmp_icb_cmd_valid_37;
  wire     tmp_icb_cmd_ready_37;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_37 (
    .i_vld(tmp_icb_cmd_valid_36), 
    .i_rdy(tmp_icb_cmd_ready_36), 
    .i_dat(tmp_icb_cmd_pack_36),
    .o_vld(tmp_icb_cmd_valid_37), 
    .o_rdy(delay_stage_select[37] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_37), 
    .o_dat(tmp_icb_cmd_pack_37),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_38;
  wire     tmp_icb_cmd_valid_38;
  wire     tmp_icb_cmd_ready_38;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_38 (
    .i_vld(tmp_icb_cmd_valid_37), 
    .i_rdy(tmp_icb_cmd_ready_37), 
    .i_dat(tmp_icb_cmd_pack_37),
    .o_vld(tmp_icb_cmd_valid_38), 
    .o_rdy(delay_stage_select[38] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_38), 
    .o_dat(tmp_icb_cmd_pack_38),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_39;
  wire     tmp_icb_cmd_valid_39;
  wire     tmp_icb_cmd_ready_39;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_39 (
    .i_vld(tmp_icb_cmd_valid_38), 
    .i_rdy(tmp_icb_cmd_ready_38), 
    .i_dat(tmp_icb_cmd_pack_38),
    .o_vld(tmp_icb_cmd_valid_39), 
    .o_rdy(delay_stage_select[39] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_39), 
    .o_dat(tmp_icb_cmd_pack_39),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_40;
  wire     tmp_icb_cmd_valid_40;
  wire     tmp_icb_cmd_ready_40;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_40 (
    .i_vld(tmp_icb_cmd_valid_39), 
    .i_rdy(tmp_icb_cmd_ready_39), 
    .i_dat(tmp_icb_cmd_pack_39),
    .o_vld(tmp_icb_cmd_valid_40), 
    .o_rdy(delay_stage_select[40] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_40), 
    .o_dat(tmp_icb_cmd_pack_40),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_41;
  wire     tmp_icb_cmd_valid_41;
  wire     tmp_icb_cmd_ready_41;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_41 (
    .i_vld(tmp_icb_cmd_valid_40), 
    .i_rdy(tmp_icb_cmd_ready_40), 
    .i_dat(tmp_icb_cmd_pack_40),
    .o_vld(tmp_icb_cmd_valid_41), 
    .o_rdy(delay_stage_select[41] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_41), 
    .o_dat(tmp_icb_cmd_pack_41),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_42;
  wire     tmp_icb_cmd_valid_42;
  wire     tmp_icb_cmd_ready_42;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_42 (
    .i_vld(tmp_icb_cmd_valid_41), 
    .i_rdy(tmp_icb_cmd_ready_41), 
    .i_dat(tmp_icb_cmd_pack_41),
    .o_vld(tmp_icb_cmd_valid_42), 
    .o_rdy(delay_stage_select[42] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_42), 
    .o_dat(tmp_icb_cmd_pack_42),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_43;
  wire     tmp_icb_cmd_valid_43;
  wire     tmp_icb_cmd_ready_43;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_43 (
    .i_vld(tmp_icb_cmd_valid_42), 
    .i_rdy(tmp_icb_cmd_ready_42), 
    .i_dat(tmp_icb_cmd_pack_42),
    .o_vld(tmp_icb_cmd_valid_43), 
    .o_rdy(delay_stage_select[43] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_43), 
    .o_dat(tmp_icb_cmd_pack_43),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_44;
  wire     tmp_icb_cmd_valid_44;
  wire     tmp_icb_cmd_ready_44;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_44 (
    .i_vld(tmp_icb_cmd_valid_43), 
    .i_rdy(tmp_icb_cmd_ready_43), 
    .i_dat(tmp_icb_cmd_pack_43),
    .o_vld(tmp_icb_cmd_valid_44), 
    .o_rdy(delay_stage_select[44] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_44), 
    .o_dat(tmp_icb_cmd_pack_44),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_45;
  wire     tmp_icb_cmd_valid_45;
  wire     tmp_icb_cmd_ready_45;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_45 (
    .i_vld(tmp_icb_cmd_valid_44), 
    .i_rdy(tmp_icb_cmd_ready_44), 
    .i_dat(tmp_icb_cmd_pack_44),
    .o_vld(tmp_icb_cmd_valid_45), 
    .o_rdy(delay_stage_select[45] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_45), 
    .o_dat(tmp_icb_cmd_pack_45),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_46;
  wire     tmp_icb_cmd_valid_46;
  wire     tmp_icb_cmd_ready_46;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_46 (
    .i_vld(tmp_icb_cmd_valid_45), 
    .i_rdy(tmp_icb_cmd_ready_45), 
    .i_dat(tmp_icb_cmd_pack_45),
    .o_vld(tmp_icb_cmd_valid_46), 
    .o_rdy(delay_stage_select[46] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_46), 
    .o_dat(tmp_icb_cmd_pack_46),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_47;
  wire     tmp_icb_cmd_valid_47;
  wire     tmp_icb_cmd_ready_47;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_47 (
    .i_vld(tmp_icb_cmd_valid_46), 
    .i_rdy(tmp_icb_cmd_ready_46), 
    .i_dat(tmp_icb_cmd_pack_46),
    .o_vld(tmp_icb_cmd_valid_47), 
    .o_rdy(delay_stage_select[47] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_47), 
    .o_dat(tmp_icb_cmd_pack_47),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_48;
  wire     tmp_icb_cmd_valid_48;
  wire     tmp_icb_cmd_ready_48;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_48 (
    .i_vld(tmp_icb_cmd_valid_47), 
    .i_rdy(tmp_icb_cmd_ready_47), 
    .i_dat(tmp_icb_cmd_pack_47),
    .o_vld(tmp_icb_cmd_valid_48), 
    .o_rdy(delay_stage_select[48] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_48), 
    .o_dat(tmp_icb_cmd_pack_48),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_49;
  wire     tmp_icb_cmd_valid_49;
  wire     tmp_icb_cmd_ready_49;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_49 (
    .i_vld(tmp_icb_cmd_valid_48), 
    .i_rdy(tmp_icb_cmd_ready_48), 
    .i_dat(tmp_icb_cmd_pack_48),
    .o_vld(tmp_icb_cmd_valid_49), 
    .o_rdy(delay_stage_select[49] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_49), 
    .o_dat(tmp_icb_cmd_pack_49),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_50;
  wire     tmp_icb_cmd_valid_50;
  wire     tmp_icb_cmd_ready_50;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_50 (
    .i_vld(tmp_icb_cmd_valid_49), 
    .i_rdy(tmp_icb_cmd_ready_49), 
    .i_dat(tmp_icb_cmd_pack_49),
    .o_vld(tmp_icb_cmd_valid_50), 
    .o_rdy(delay_stage_select[50] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_50), 
    .o_dat(tmp_icb_cmd_pack_50),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_51;
  wire     tmp_icb_cmd_valid_51;
  wire     tmp_icb_cmd_ready_51;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_51 (
    .i_vld(tmp_icb_cmd_valid_50), 
    .i_rdy(tmp_icb_cmd_ready_50), 
    .i_dat(tmp_icb_cmd_pack_50),
    .o_vld(tmp_icb_cmd_valid_51), 
    .o_rdy(delay_stage_select[51] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_51), 
    .o_dat(tmp_icb_cmd_pack_51),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_52;
  wire     tmp_icb_cmd_valid_52;
  wire     tmp_icb_cmd_ready_52;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_52 (
    .i_vld(tmp_icb_cmd_valid_51), 
    .i_rdy(tmp_icb_cmd_ready_51), 
    .i_dat(tmp_icb_cmd_pack_51),
    .o_vld(tmp_icb_cmd_valid_52), 
    .o_rdy(delay_stage_select[52] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_52), 
    .o_dat(tmp_icb_cmd_pack_52),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_53;
  wire     tmp_icb_cmd_valid_53;
  wire     tmp_icb_cmd_ready_53;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_53 (
    .i_vld(tmp_icb_cmd_valid_52), 
    .i_rdy(tmp_icb_cmd_ready_52), 
    .i_dat(tmp_icb_cmd_pack_52),
    .o_vld(tmp_icb_cmd_valid_53), 
    .o_rdy(delay_stage_select[53] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_53), 
    .o_dat(tmp_icb_cmd_pack_53),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_54;
  wire     tmp_icb_cmd_valid_54;
  wire     tmp_icb_cmd_ready_54;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_54 (
    .i_vld(tmp_icb_cmd_valid_53), 
    .i_rdy(tmp_icb_cmd_ready_53), 
    .i_dat(tmp_icb_cmd_pack_53),
    .o_vld(tmp_icb_cmd_valid_54), 
    .o_rdy(delay_stage_select[54] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_54), 
    .o_dat(tmp_icb_cmd_pack_54),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_55;
  wire     tmp_icb_cmd_valid_55;
  wire     tmp_icb_cmd_ready_55;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_55 (
    .i_vld(tmp_icb_cmd_valid_54), 
    .i_rdy(tmp_icb_cmd_ready_54), 
    .i_dat(tmp_icb_cmd_pack_54),
    .o_vld(tmp_icb_cmd_valid_55), 
    .o_rdy(delay_stage_select[55] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_55), 
    .o_dat(tmp_icb_cmd_pack_55),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_56;
  wire     tmp_icb_cmd_valid_56;
  wire     tmp_icb_cmd_ready_56;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_56 (
    .i_vld(tmp_icb_cmd_valid_55), 
    .i_rdy(tmp_icb_cmd_ready_55), 
    .i_dat(tmp_icb_cmd_pack_55),
    .o_vld(tmp_icb_cmd_valid_56), 
    .o_rdy(delay_stage_select[56] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_56), 
    .o_dat(tmp_icb_cmd_pack_56),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_57;
  wire     tmp_icb_cmd_valid_57;
  wire     tmp_icb_cmd_ready_57;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_57 (
    .i_vld(tmp_icb_cmd_valid_56), 
    .i_rdy(tmp_icb_cmd_ready_56), 
    .i_dat(tmp_icb_cmd_pack_56),
    .o_vld(tmp_icb_cmd_valid_57), 
    .o_rdy(delay_stage_select[57] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_57), 
    .o_dat(tmp_icb_cmd_pack_57),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_58;
  wire     tmp_icb_cmd_valid_58;
  wire     tmp_icb_cmd_ready_58;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_58 (
    .i_vld(tmp_icb_cmd_valid_57), 
    .i_rdy(tmp_icb_cmd_ready_57), 
    .i_dat(tmp_icb_cmd_pack_57),
    .o_vld(tmp_icb_cmd_valid_58), 
    .o_rdy(delay_stage_select[58] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_58), 
    .o_dat(tmp_icb_cmd_pack_58),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_59;
  wire     tmp_icb_cmd_valid_59;
  wire     tmp_icb_cmd_ready_59;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_59 (
    .i_vld(tmp_icb_cmd_valid_58), 
    .i_rdy(tmp_icb_cmd_ready_58), 
    .i_dat(tmp_icb_cmd_pack_58),
    .o_vld(tmp_icb_cmd_valid_59), 
    .o_rdy(delay_stage_select[59] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_59), 
    .o_dat(tmp_icb_cmd_pack_59),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_60;
  wire     tmp_icb_cmd_valid_60;
  wire     tmp_icb_cmd_ready_60;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_60 (
    .i_vld(tmp_icb_cmd_valid_59), 
    .i_rdy(tmp_icb_cmd_ready_59), 
    .i_dat(tmp_icb_cmd_pack_59),
    .o_vld(tmp_icb_cmd_valid_60), 
    .o_rdy(delay_stage_select[60] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_60), 
    .o_dat(tmp_icb_cmd_pack_60),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_61;
  wire     tmp_icb_cmd_valid_61;
  wire     tmp_icb_cmd_ready_61;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_61 (
    .i_vld(tmp_icb_cmd_valid_60), 
    .i_rdy(tmp_icb_cmd_ready_60), 
    .i_dat(tmp_icb_cmd_pack_60),
    .o_vld(tmp_icb_cmd_valid_61), 
    .o_rdy(delay_stage_select[61] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_61), 
    .o_dat(tmp_icb_cmd_pack_61),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_62;
  wire     tmp_icb_cmd_valid_62;
  wire     tmp_icb_cmd_ready_62;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_62 (
    .i_vld(tmp_icb_cmd_valid_61), 
    .i_rdy(tmp_icb_cmd_ready_61), 
    .i_dat(tmp_icb_cmd_pack_61),
    .o_vld(tmp_icb_cmd_valid_62), 
    .o_rdy(delay_stage_select[62] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_62), 
    .o_dat(tmp_icb_cmd_pack_62),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_63;
  wire     tmp_icb_cmd_valid_63;
  wire     tmp_icb_cmd_ready_63;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_63 (
    .i_vld(tmp_icb_cmd_valid_62), 
    .i_rdy(tmp_icb_cmd_ready_62), 
    .i_dat(tmp_icb_cmd_pack_62),
    .o_vld(tmp_icb_cmd_valid_63), 
    .o_rdy(delay_stage_select[63] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_63), 
    .o_dat(tmp_icb_cmd_pack_63),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_64;
  wire     tmp_icb_cmd_valid_64;
  wire     tmp_icb_cmd_ready_64;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_64 (
    .i_vld(tmp_icb_cmd_valid_63), 
    .i_rdy(tmp_icb_cmd_ready_63), 
    .i_dat(tmp_icb_cmd_pack_63),
    .o_vld(tmp_icb_cmd_valid_64), 
    .o_rdy(delay_stage_select[64] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_64), 
    .o_dat(tmp_icb_cmd_pack_64),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_65;
  wire     tmp_icb_cmd_valid_65;
  wire     tmp_icb_cmd_ready_65;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_65 (
    .i_vld(tmp_icb_cmd_valid_64), 
    .i_rdy(tmp_icb_cmd_ready_64), 
    .i_dat(tmp_icb_cmd_pack_64),
    .o_vld(tmp_icb_cmd_valid_65), 
    .o_rdy(delay_stage_select[65] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_65), 
    .o_dat(tmp_icb_cmd_pack_65),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_66;
  wire     tmp_icb_cmd_valid_66;
  wire     tmp_icb_cmd_ready_66;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_66 (
    .i_vld(tmp_icb_cmd_valid_65), 
    .i_rdy(tmp_icb_cmd_ready_65), 
    .i_dat(tmp_icb_cmd_pack_65),
    .o_vld(tmp_icb_cmd_valid_66), 
    .o_rdy(delay_stage_select[66] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_66), 
    .o_dat(tmp_icb_cmd_pack_66),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_67;
  wire     tmp_icb_cmd_valid_67;
  wire     tmp_icb_cmd_ready_67;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_67 (
    .i_vld(tmp_icb_cmd_valid_66), 
    .i_rdy(tmp_icb_cmd_ready_66), 
    .i_dat(tmp_icb_cmd_pack_66),
    .o_vld(tmp_icb_cmd_valid_67), 
    .o_rdy(delay_stage_select[67] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_67), 
    .o_dat(tmp_icb_cmd_pack_67),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_68;
  wire     tmp_icb_cmd_valid_68;
  wire     tmp_icb_cmd_ready_68;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_68 (
    .i_vld(tmp_icb_cmd_valid_67), 
    .i_rdy(tmp_icb_cmd_ready_67), 
    .i_dat(tmp_icb_cmd_pack_67),
    .o_vld(tmp_icb_cmd_valid_68), 
    .o_rdy(delay_stage_select[68] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_68), 
    .o_dat(tmp_icb_cmd_pack_68),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_69;
  wire     tmp_icb_cmd_valid_69;
  wire     tmp_icb_cmd_ready_69;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_69 (
    .i_vld(tmp_icb_cmd_valid_68), 
    .i_rdy(tmp_icb_cmd_ready_68), 
    .i_dat(tmp_icb_cmd_pack_68),
    .o_vld(tmp_icb_cmd_valid_69), 
    .o_rdy(delay_stage_select[69] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_69), 
    .o_dat(tmp_icb_cmd_pack_69),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_70;
  wire     tmp_icb_cmd_valid_70;
  wire     tmp_icb_cmd_ready_70;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_70 (
    .i_vld(tmp_icb_cmd_valid_69), 
    .i_rdy(tmp_icb_cmd_ready_69), 
    .i_dat(tmp_icb_cmd_pack_69),
    .o_vld(tmp_icb_cmd_valid_70), 
    .o_rdy(delay_stage_select[70] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_70), 
    .o_dat(tmp_icb_cmd_pack_70),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_71;
  wire     tmp_icb_cmd_valid_71;
  wire     tmp_icb_cmd_ready_71;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_71 (
    .i_vld(tmp_icb_cmd_valid_70), 
    .i_rdy(tmp_icb_cmd_ready_70), 
    .i_dat(tmp_icb_cmd_pack_70),
    .o_vld(tmp_icb_cmd_valid_71), 
    .o_rdy(delay_stage_select[71] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_71), 
    .o_dat(tmp_icb_cmd_pack_71),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_72;
  wire     tmp_icb_cmd_valid_72;
  wire     tmp_icb_cmd_ready_72;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_72 (
    .i_vld(tmp_icb_cmd_valid_71), 
    .i_rdy(tmp_icb_cmd_ready_71), 
    .i_dat(tmp_icb_cmd_pack_71),
    .o_vld(tmp_icb_cmd_valid_72), 
    .o_rdy(delay_stage_select[72] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_72), 
    .o_dat(tmp_icb_cmd_pack_72),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_73;
  wire     tmp_icb_cmd_valid_73;
  wire     tmp_icb_cmd_ready_73;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_73 (
    .i_vld(tmp_icb_cmd_valid_72), 
    .i_rdy(tmp_icb_cmd_ready_72), 
    .i_dat(tmp_icb_cmd_pack_72),
    .o_vld(tmp_icb_cmd_valid_73), 
    .o_rdy(delay_stage_select[73] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_73), 
    .o_dat(tmp_icb_cmd_pack_73),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_74;
  wire     tmp_icb_cmd_valid_74;
  wire     tmp_icb_cmd_ready_74;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_74 (
    .i_vld(tmp_icb_cmd_valid_73), 
    .i_rdy(tmp_icb_cmd_ready_73), 
    .i_dat(tmp_icb_cmd_pack_73),
    .o_vld(tmp_icb_cmd_valid_74), 
    .o_rdy(delay_stage_select[74] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_74), 
    .o_dat(tmp_icb_cmd_pack_74),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_75;
  wire     tmp_icb_cmd_valid_75;
  wire     tmp_icb_cmd_ready_75;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_75 (
    .i_vld(tmp_icb_cmd_valid_74), 
    .i_rdy(tmp_icb_cmd_ready_74), 
    .i_dat(tmp_icb_cmd_pack_74),
    .o_vld(tmp_icb_cmd_valid_75), 
    .o_rdy(delay_stage_select[75] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_75), 
    .o_dat(tmp_icb_cmd_pack_75),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_76;
  wire     tmp_icb_cmd_valid_76;
  wire     tmp_icb_cmd_ready_76;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_76 (
    .i_vld(tmp_icb_cmd_valid_75), 
    .i_rdy(tmp_icb_cmd_ready_75), 
    .i_dat(tmp_icb_cmd_pack_75),
    .o_vld(tmp_icb_cmd_valid_76), 
    .o_rdy(delay_stage_select[76] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_76), 
    .o_dat(tmp_icb_cmd_pack_76),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_77;
  wire     tmp_icb_cmd_valid_77;
  wire     tmp_icb_cmd_ready_77;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_77 (
    .i_vld(tmp_icb_cmd_valid_76), 
    .i_rdy(tmp_icb_cmd_ready_76), 
    .i_dat(tmp_icb_cmd_pack_76),
    .o_vld(tmp_icb_cmd_valid_77), 
    .o_rdy(delay_stage_select[77] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_77), 
    .o_dat(tmp_icb_cmd_pack_77),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_78;
  wire     tmp_icb_cmd_valid_78;
  wire     tmp_icb_cmd_ready_78;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_78 (
    .i_vld(tmp_icb_cmd_valid_77), 
    .i_rdy(tmp_icb_cmd_ready_77), 
    .i_dat(tmp_icb_cmd_pack_77),
    .o_vld(tmp_icb_cmd_valid_78), 
    .o_rdy(delay_stage_select[78] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_78), 
    .o_dat(tmp_icb_cmd_pack_78),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_79;
  wire     tmp_icb_cmd_valid_79;
  wire     tmp_icb_cmd_ready_79;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_79 (
    .i_vld(tmp_icb_cmd_valid_78), 
    .i_rdy(tmp_icb_cmd_ready_78), 
    .i_dat(tmp_icb_cmd_pack_78),
    .o_vld(tmp_icb_cmd_valid_79), 
    .o_rdy(delay_stage_select[79] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_79), 
    .o_dat(tmp_icb_cmd_pack_79),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_80;
  wire     tmp_icb_cmd_valid_80;
  wire     tmp_icb_cmd_ready_80;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_80 (
    .i_vld(tmp_icb_cmd_valid_79), 
    .i_rdy(tmp_icb_cmd_ready_79), 
    .i_dat(tmp_icb_cmd_pack_79),
    .o_vld(tmp_icb_cmd_valid_80), 
    .o_rdy(delay_stage_select[80] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_80), 
    .o_dat(tmp_icb_cmd_pack_80),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_81;
  wire     tmp_icb_cmd_valid_81;
  wire     tmp_icb_cmd_ready_81;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_81 (
    .i_vld(tmp_icb_cmd_valid_80), 
    .i_rdy(tmp_icb_cmd_ready_80), 
    .i_dat(tmp_icb_cmd_pack_80),
    .o_vld(tmp_icb_cmd_valid_81), 
    .o_rdy(delay_stage_select[81] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_81), 
    .o_dat(tmp_icb_cmd_pack_81),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_82;
  wire     tmp_icb_cmd_valid_82;
  wire     tmp_icb_cmd_ready_82;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_82 (
    .i_vld(tmp_icb_cmd_valid_81), 
    .i_rdy(tmp_icb_cmd_ready_81), 
    .i_dat(tmp_icb_cmd_pack_81),
    .o_vld(tmp_icb_cmd_valid_82), 
    .o_rdy(delay_stage_select[82] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_82), 
    .o_dat(tmp_icb_cmd_pack_82),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_83;
  wire     tmp_icb_cmd_valid_83;
  wire     tmp_icb_cmd_ready_83;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_83 (
    .i_vld(tmp_icb_cmd_valid_82), 
    .i_rdy(tmp_icb_cmd_ready_82), 
    .i_dat(tmp_icb_cmd_pack_82),
    .o_vld(tmp_icb_cmd_valid_83), 
    .o_rdy(delay_stage_select[83] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_83), 
    .o_dat(tmp_icb_cmd_pack_83),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_84;
  wire     tmp_icb_cmd_valid_84;
  wire     tmp_icb_cmd_ready_84;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_84 (
    .i_vld(tmp_icb_cmd_valid_83), 
    .i_rdy(tmp_icb_cmd_ready_83), 
    .i_dat(tmp_icb_cmd_pack_83),
    .o_vld(tmp_icb_cmd_valid_84), 
    .o_rdy(delay_stage_select[84] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_84), 
    .o_dat(tmp_icb_cmd_pack_84),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_85;
  wire     tmp_icb_cmd_valid_85;
  wire     tmp_icb_cmd_ready_85;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_85 (
    .i_vld(tmp_icb_cmd_valid_84), 
    .i_rdy(tmp_icb_cmd_ready_84), 
    .i_dat(tmp_icb_cmd_pack_84),
    .o_vld(tmp_icb_cmd_valid_85), 
    .o_rdy(delay_stage_select[85] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_85), 
    .o_dat(tmp_icb_cmd_pack_85),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_86;
  wire     tmp_icb_cmd_valid_86;
  wire     tmp_icb_cmd_ready_86;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_86 (
    .i_vld(tmp_icb_cmd_valid_85), 
    .i_rdy(tmp_icb_cmd_ready_85), 
    .i_dat(tmp_icb_cmd_pack_85),
    .o_vld(tmp_icb_cmd_valid_86), 
    .o_rdy(delay_stage_select[86] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_86), 
    .o_dat(tmp_icb_cmd_pack_86),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_87;
  wire     tmp_icb_cmd_valid_87;
  wire     tmp_icb_cmd_ready_87;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_87 (
    .i_vld(tmp_icb_cmd_valid_86), 
    .i_rdy(tmp_icb_cmd_ready_86), 
    .i_dat(tmp_icb_cmd_pack_86),
    .o_vld(tmp_icb_cmd_valid_87), 
    .o_rdy(delay_stage_select[87] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_87), 
    .o_dat(tmp_icb_cmd_pack_87),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_88;
  wire     tmp_icb_cmd_valid_88;
  wire     tmp_icb_cmd_ready_88;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_88 (
    .i_vld(tmp_icb_cmd_valid_87), 
    .i_rdy(tmp_icb_cmd_ready_87), 
    .i_dat(tmp_icb_cmd_pack_87),
    .o_vld(tmp_icb_cmd_valid_88), 
    .o_rdy(delay_stage_select[88] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_88), 
    .o_dat(tmp_icb_cmd_pack_88),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_89;
  wire     tmp_icb_cmd_valid_89;
  wire     tmp_icb_cmd_ready_89;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_89 (
    .i_vld(tmp_icb_cmd_valid_88), 
    .i_rdy(tmp_icb_cmd_ready_88), 
    .i_dat(tmp_icb_cmd_pack_88),
    .o_vld(tmp_icb_cmd_valid_89), 
    .o_rdy(delay_stage_select[89] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_89), 
    .o_dat(tmp_icb_cmd_pack_89),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_90;
  wire     tmp_icb_cmd_valid_90;
  wire     tmp_icb_cmd_ready_90;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_90 (
    .i_vld(tmp_icb_cmd_valid_89), 
    .i_rdy(tmp_icb_cmd_ready_89), 
    .i_dat(tmp_icb_cmd_pack_89),
    .o_vld(tmp_icb_cmd_valid_90), 
    .o_rdy(delay_stage_select[90] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_90), 
    .o_dat(tmp_icb_cmd_pack_90),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_91;
  wire     tmp_icb_cmd_valid_91;
  wire     tmp_icb_cmd_ready_91;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_91 (
    .i_vld(tmp_icb_cmd_valid_90), 
    .i_rdy(tmp_icb_cmd_ready_90), 
    .i_dat(tmp_icb_cmd_pack_90),
    .o_vld(tmp_icb_cmd_valid_91), 
    .o_rdy(delay_stage_select[91] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_91), 
    .o_dat(tmp_icb_cmd_pack_91),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_92;
  wire     tmp_icb_cmd_valid_92;
  wire     tmp_icb_cmd_ready_92;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_92 (
    .i_vld(tmp_icb_cmd_valid_91), 
    .i_rdy(tmp_icb_cmd_ready_91), 
    .i_dat(tmp_icb_cmd_pack_91),
    .o_vld(tmp_icb_cmd_valid_92), 
    .o_rdy(delay_stage_select[92] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_92), 
    .o_dat(tmp_icb_cmd_pack_92),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_93;
  wire     tmp_icb_cmd_valid_93;
  wire     tmp_icb_cmd_ready_93;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_93 (
    .i_vld(tmp_icb_cmd_valid_92), 
    .i_rdy(tmp_icb_cmd_ready_92), 
    .i_dat(tmp_icb_cmd_pack_92),
    .o_vld(tmp_icb_cmd_valid_93), 
    .o_rdy(delay_stage_select[93] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_93), 
    .o_dat(tmp_icb_cmd_pack_93),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_94;
  wire     tmp_icb_cmd_valid_94;
  wire     tmp_icb_cmd_ready_94;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_94 (
    .i_vld(tmp_icb_cmd_valid_93), 
    .i_rdy(tmp_icb_cmd_ready_93), 
    .i_dat(tmp_icb_cmd_pack_93),
    .o_vld(tmp_icb_cmd_valid_94), 
    .o_rdy(delay_stage_select[94] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_94), 
    .o_dat(tmp_icb_cmd_pack_94),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_95;
  wire     tmp_icb_cmd_valid_95;
  wire     tmp_icb_cmd_ready_95;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_95 (
    .i_vld(tmp_icb_cmd_valid_94), 
    .i_rdy(tmp_icb_cmd_ready_94), 
    .i_dat(tmp_icb_cmd_pack_94),
    .o_vld(tmp_icb_cmd_valid_95), 
    .o_rdy(delay_stage_select[95] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_95), 
    .o_dat(tmp_icb_cmd_pack_95),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_96;
  wire     tmp_icb_cmd_valid_96;
  wire     tmp_icb_cmd_ready_96;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_96 (
    .i_vld(tmp_icb_cmd_valid_95), 
    .i_rdy(tmp_icb_cmd_ready_95), 
    .i_dat(tmp_icb_cmd_pack_95),
    .o_vld(tmp_icb_cmd_valid_96), 
    .o_rdy(delay_stage_select[96] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_96), 
    .o_dat(tmp_icb_cmd_pack_96),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_97;
  wire     tmp_icb_cmd_valid_97;
  wire     tmp_icb_cmd_ready_97;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_97 (
    .i_vld(tmp_icb_cmd_valid_96), 
    .i_rdy(tmp_icb_cmd_ready_96), 
    .i_dat(tmp_icb_cmd_pack_96),
    .o_vld(tmp_icb_cmd_valid_97), 
    .o_rdy(delay_stage_select[97] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_97), 
    .o_dat(tmp_icb_cmd_pack_97),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_98;
  wire     tmp_icb_cmd_valid_98;
  wire     tmp_icb_cmd_ready_98;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_98 (
    .i_vld(tmp_icb_cmd_valid_97), 
    .i_rdy(tmp_icb_cmd_ready_97), 
    .i_dat(tmp_icb_cmd_pack_97),
    .o_vld(tmp_icb_cmd_valid_98), 
    .o_rdy(delay_stage_select[98] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_98), 
    .o_dat(tmp_icb_cmd_pack_98),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_99;
  wire     tmp_icb_cmd_valid_99;
  wire     tmp_icb_cmd_ready_99;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_99 (
    .i_vld(tmp_icb_cmd_valid_98), 
    .i_rdy(tmp_icb_cmd_ready_98), 
    .i_dat(tmp_icb_cmd_pack_98),
    .o_vld(tmp_icb_cmd_valid_99), 
    .o_rdy(delay_stage_select[99] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_99), 
    .o_dat(tmp_icb_cmd_pack_99),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_100;
  wire     tmp_icb_cmd_valid_100;
  wire     tmp_icb_cmd_ready_100;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_100 (
    .i_vld(tmp_icb_cmd_valid_99), 
    .i_rdy(tmp_icb_cmd_ready_99), 
    .i_dat(tmp_icb_cmd_pack_99),
    .o_vld(tmp_icb_cmd_valid_100), 
    .o_rdy(delay_stage_select[100] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_100), 
    .o_dat(tmp_icb_cmd_pack_100),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_101;
  wire     tmp_icb_cmd_valid_101;
  wire     tmp_icb_cmd_ready_101;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_101 (
    .i_vld(tmp_icb_cmd_valid_100), 
    .i_rdy(tmp_icb_cmd_ready_100), 
    .i_dat(tmp_icb_cmd_pack_100),
    .o_vld(tmp_icb_cmd_valid_101), 
    .o_rdy(delay_stage_select[101] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_101), 
    .o_dat(tmp_icb_cmd_pack_101),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_102;
  wire     tmp_icb_cmd_valid_102;
  wire     tmp_icb_cmd_ready_102;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_102 (
    .i_vld(tmp_icb_cmd_valid_101), 
    .i_rdy(tmp_icb_cmd_ready_101), 
    .i_dat(tmp_icb_cmd_pack_101),
    .o_vld(tmp_icb_cmd_valid_102), 
    .o_rdy(delay_stage_select[102] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_102), 
    .o_dat(tmp_icb_cmd_pack_102),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_103;
  wire     tmp_icb_cmd_valid_103;
  wire     tmp_icb_cmd_ready_103;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_103 (
    .i_vld(tmp_icb_cmd_valid_102), 
    .i_rdy(tmp_icb_cmd_ready_102), 
    .i_dat(tmp_icb_cmd_pack_102),
    .o_vld(tmp_icb_cmd_valid_103), 
    .o_rdy(delay_stage_select[103] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_103), 
    .o_dat(tmp_icb_cmd_pack_103),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_104;
  wire     tmp_icb_cmd_valid_104;
  wire     tmp_icb_cmd_ready_104;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_104 (
    .i_vld(tmp_icb_cmd_valid_103), 
    .i_rdy(tmp_icb_cmd_ready_103), 
    .i_dat(tmp_icb_cmd_pack_103),
    .o_vld(tmp_icb_cmd_valid_104), 
    .o_rdy(delay_stage_select[104] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_104), 
    .o_dat(tmp_icb_cmd_pack_104),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_105;
  wire     tmp_icb_cmd_valid_105;
  wire     tmp_icb_cmd_ready_105;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_105 (
    .i_vld(tmp_icb_cmd_valid_104), 
    .i_rdy(tmp_icb_cmd_ready_104), 
    .i_dat(tmp_icb_cmd_pack_104),
    .o_vld(tmp_icb_cmd_valid_105), 
    .o_rdy(delay_stage_select[105] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_105), 
    .o_dat(tmp_icb_cmd_pack_105),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_106;
  wire     tmp_icb_cmd_valid_106;
  wire     tmp_icb_cmd_ready_106;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_106 (
    .i_vld(tmp_icb_cmd_valid_105), 
    .i_rdy(tmp_icb_cmd_ready_105), 
    .i_dat(tmp_icb_cmd_pack_105),
    .o_vld(tmp_icb_cmd_valid_106), 
    .o_rdy(delay_stage_select[106] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_106), 
    .o_dat(tmp_icb_cmd_pack_106),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_107;
  wire     tmp_icb_cmd_valid_107;
  wire     tmp_icb_cmd_ready_107;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_107 (
    .i_vld(tmp_icb_cmd_valid_106), 
    .i_rdy(tmp_icb_cmd_ready_106), 
    .i_dat(tmp_icb_cmd_pack_106),
    .o_vld(tmp_icb_cmd_valid_107), 
    .o_rdy(delay_stage_select[107] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_107), 
    .o_dat(tmp_icb_cmd_pack_107),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_108;
  wire     tmp_icb_cmd_valid_108;
  wire     tmp_icb_cmd_ready_108;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_108 (
    .i_vld(tmp_icb_cmd_valid_107), 
    .i_rdy(tmp_icb_cmd_ready_107), 
    .i_dat(tmp_icb_cmd_pack_107),
    .o_vld(tmp_icb_cmd_valid_108), 
    .o_rdy(delay_stage_select[108] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_108), 
    .o_dat(tmp_icb_cmd_pack_108),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_109;
  wire     tmp_icb_cmd_valid_109;
  wire     tmp_icb_cmd_ready_109;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_109 (
    .i_vld(tmp_icb_cmd_valid_108), 
    .i_rdy(tmp_icb_cmd_ready_108), 
    .i_dat(tmp_icb_cmd_pack_108),
    .o_vld(tmp_icb_cmd_valid_109), 
    .o_rdy(delay_stage_select[109] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_109), 
    .o_dat(tmp_icb_cmd_pack_109),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_110;
  wire     tmp_icb_cmd_valid_110;
  wire     tmp_icb_cmd_ready_110;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_110 (
    .i_vld(tmp_icb_cmd_valid_109), 
    .i_rdy(tmp_icb_cmd_ready_109), 
    .i_dat(tmp_icb_cmd_pack_109),
    .o_vld(tmp_icb_cmd_valid_110), 
    .o_rdy(delay_stage_select[110] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_110), 
    .o_dat(tmp_icb_cmd_pack_110),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_111;
  wire     tmp_icb_cmd_valid_111;
  wire     tmp_icb_cmd_ready_111;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_111 (
    .i_vld(tmp_icb_cmd_valid_110), 
    .i_rdy(tmp_icb_cmd_ready_110), 
    .i_dat(tmp_icb_cmd_pack_110),
    .o_vld(tmp_icb_cmd_valid_111), 
    .o_rdy(delay_stage_select[111] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_111), 
    .o_dat(tmp_icb_cmd_pack_111),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_112;
  wire     tmp_icb_cmd_valid_112;
  wire     tmp_icb_cmd_ready_112;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_112 (
    .i_vld(tmp_icb_cmd_valid_111), 
    .i_rdy(tmp_icb_cmd_ready_111), 
    .i_dat(tmp_icb_cmd_pack_111),
    .o_vld(tmp_icb_cmd_valid_112), 
    .o_rdy(delay_stage_select[112] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_112), 
    .o_dat(tmp_icb_cmd_pack_112),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_113;
  wire     tmp_icb_cmd_valid_113;
  wire     tmp_icb_cmd_ready_113;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_113 (
    .i_vld(tmp_icb_cmd_valid_112), 
    .i_rdy(tmp_icb_cmd_ready_112), 
    .i_dat(tmp_icb_cmd_pack_112),
    .o_vld(tmp_icb_cmd_valid_113), 
    .o_rdy(delay_stage_select[113] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_113), 
    .o_dat(tmp_icb_cmd_pack_113),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_114;
  wire     tmp_icb_cmd_valid_114;
  wire     tmp_icb_cmd_ready_114;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_114 (
    .i_vld(tmp_icb_cmd_valid_113), 
    .i_rdy(tmp_icb_cmd_ready_113), 
    .i_dat(tmp_icb_cmd_pack_113),
    .o_vld(tmp_icb_cmd_valid_114), 
    .o_rdy(delay_stage_select[114] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_114), 
    .o_dat(tmp_icb_cmd_pack_114),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_115;
  wire     tmp_icb_cmd_valid_115;
  wire     tmp_icb_cmd_ready_115;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_115 (
    .i_vld(tmp_icb_cmd_valid_114), 
    .i_rdy(tmp_icb_cmd_ready_114), 
    .i_dat(tmp_icb_cmd_pack_114),
    .o_vld(tmp_icb_cmd_valid_115), 
    .o_rdy(delay_stage_select[115] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_115), 
    .o_dat(tmp_icb_cmd_pack_115),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_116;
  wire     tmp_icb_cmd_valid_116;
  wire     tmp_icb_cmd_ready_116;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_116 (
    .i_vld(tmp_icb_cmd_valid_115), 
    .i_rdy(tmp_icb_cmd_ready_115), 
    .i_dat(tmp_icb_cmd_pack_115),
    .o_vld(tmp_icb_cmd_valid_116), 
    .o_rdy(delay_stage_select[116] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_116), 
    .o_dat(tmp_icb_cmd_pack_116),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_117;
  wire     tmp_icb_cmd_valid_117;
  wire     tmp_icb_cmd_ready_117;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_117 (
    .i_vld(tmp_icb_cmd_valid_116), 
    .i_rdy(tmp_icb_cmd_ready_116), 
    .i_dat(tmp_icb_cmd_pack_116),
    .o_vld(tmp_icb_cmd_valid_117), 
    .o_rdy(delay_stage_select[117] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_117), 
    .o_dat(tmp_icb_cmd_pack_117),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_118;
  wire     tmp_icb_cmd_valid_118;
  wire     tmp_icb_cmd_ready_118;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_118 (
    .i_vld(tmp_icb_cmd_valid_117), 
    .i_rdy(tmp_icb_cmd_ready_117), 
    .i_dat(tmp_icb_cmd_pack_117),
    .o_vld(tmp_icb_cmd_valid_118), 
    .o_rdy(delay_stage_select[118] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_118), 
    .o_dat(tmp_icb_cmd_pack_118),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_119;
  wire     tmp_icb_cmd_valid_119;
  wire     tmp_icb_cmd_ready_119;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_119 (
    .i_vld(tmp_icb_cmd_valid_118), 
    .i_rdy(tmp_icb_cmd_ready_118), 
    .i_dat(tmp_icb_cmd_pack_118),
    .o_vld(tmp_icb_cmd_valid_119), 
    .o_rdy(delay_stage_select[119] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_119), 
    .o_dat(tmp_icb_cmd_pack_119),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_120;
  wire     tmp_icb_cmd_valid_120;
  wire     tmp_icb_cmd_ready_120;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_120 (
    .i_vld(tmp_icb_cmd_valid_119), 
    .i_rdy(tmp_icb_cmd_ready_119), 
    .i_dat(tmp_icb_cmd_pack_119),
    .o_vld(tmp_icb_cmd_valid_120), 
    .o_rdy(delay_stage_select[120] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_120), 
    .o_dat(tmp_icb_cmd_pack_120),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_121;
  wire     tmp_icb_cmd_valid_121;
  wire     tmp_icb_cmd_ready_121;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_121 (
    .i_vld(tmp_icb_cmd_valid_120), 
    .i_rdy(tmp_icb_cmd_ready_120), 
    .i_dat(tmp_icb_cmd_pack_120),
    .o_vld(tmp_icb_cmd_valid_121), 
    .o_rdy(delay_stage_select[121] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_121), 
    .o_dat(tmp_icb_cmd_pack_121),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_122;
  wire     tmp_icb_cmd_valid_122;
  wire     tmp_icb_cmd_ready_122;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_122 (
    .i_vld(tmp_icb_cmd_valid_121), 
    .i_rdy(tmp_icb_cmd_ready_121), 
    .i_dat(tmp_icb_cmd_pack_121),
    .o_vld(tmp_icb_cmd_valid_122), 
    .o_rdy(delay_stage_select[122] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_122), 
    .o_dat(tmp_icb_cmd_pack_122),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_123;
  wire     tmp_icb_cmd_valid_123;
  wire     tmp_icb_cmd_ready_123;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_123 (
    .i_vld(tmp_icb_cmd_valid_122), 
    .i_rdy(tmp_icb_cmd_ready_122), 
    .i_dat(tmp_icb_cmd_pack_122),
    .o_vld(tmp_icb_cmd_valid_123), 
    .o_rdy(delay_stage_select[123] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_123), 
    .o_dat(tmp_icb_cmd_pack_123),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_124;
  wire     tmp_icb_cmd_valid_124;
  wire     tmp_icb_cmd_ready_124;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_124 (
    .i_vld(tmp_icb_cmd_valid_123), 
    .i_rdy(tmp_icb_cmd_ready_123), 
    .i_dat(tmp_icb_cmd_pack_123),
    .o_vld(tmp_icb_cmd_valid_124), 
    .o_rdy(delay_stage_select[124] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_124), 
    .o_dat(tmp_icb_cmd_pack_124),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_125;
  wire     tmp_icb_cmd_valid_125;
  wire     tmp_icb_cmd_ready_125;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_125 (
    .i_vld(tmp_icb_cmd_valid_124), 
    .i_rdy(tmp_icb_cmd_ready_124), 
    .i_dat(tmp_icb_cmd_pack_124),
    .o_vld(tmp_icb_cmd_valid_125), 
    .o_rdy(delay_stage_select[125] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_125), 
    .o_dat(tmp_icb_cmd_pack_125),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_126;
  wire     tmp_icb_cmd_valid_126;
  wire     tmp_icb_cmd_ready_126;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_126 (
    .i_vld(tmp_icb_cmd_valid_125), 
    .i_rdy(tmp_icb_cmd_ready_125), 
    .i_dat(tmp_icb_cmd_pack_125),
    .o_vld(tmp_icb_cmd_valid_126), 
    .o_rdy(delay_stage_select[126] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_126), 
    .o_dat(tmp_icb_cmd_pack_126),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_127;
  wire     tmp_icb_cmd_valid_127;
  wire     tmp_icb_cmd_ready_127;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_127 (
    .i_vld(tmp_icb_cmd_valid_126), 
    .i_rdy(tmp_icb_cmd_ready_126), 
    .i_dat(tmp_icb_cmd_pack_126),
    .o_vld(tmp_icb_cmd_valid_127), 
    .o_rdy(delay_stage_select[127] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_127), 
    .o_dat(tmp_icb_cmd_pack_127),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_128;
  wire     tmp_icb_cmd_valid_128;
  wire     tmp_icb_cmd_ready_128;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_128 (
    .i_vld(tmp_icb_cmd_valid_127), 
    .i_rdy(tmp_icb_cmd_ready_127), 
    .i_dat(tmp_icb_cmd_pack_127),
    .o_vld(tmp_icb_cmd_valid_128), 
    .o_rdy(delay_stage_select[128] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_128), 
    .o_dat(tmp_icb_cmd_pack_128),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_129;
  wire     tmp_icb_cmd_valid_129;
  wire     tmp_icb_cmd_ready_129;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_129 (
    .i_vld(tmp_icb_cmd_valid_128), 
    .i_rdy(tmp_icb_cmd_ready_128), 
    .i_dat(tmp_icb_cmd_pack_128),
    .o_vld(tmp_icb_cmd_valid_129), 
    .o_rdy(delay_stage_select[129] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_129), 
    .o_dat(tmp_icb_cmd_pack_129),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_130;
  wire     tmp_icb_cmd_valid_130;
  wire     tmp_icb_cmd_ready_130;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_130 (
    .i_vld(tmp_icb_cmd_valid_129), 
    .i_rdy(tmp_icb_cmd_ready_129), 
    .i_dat(tmp_icb_cmd_pack_129),
    .o_vld(tmp_icb_cmd_valid_130), 
    .o_rdy(delay_stage_select[130] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_130), 
    .o_dat(tmp_icb_cmd_pack_130),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_131;
  wire     tmp_icb_cmd_valid_131;
  wire     tmp_icb_cmd_ready_131;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_131 (
    .i_vld(tmp_icb_cmd_valid_130), 
    .i_rdy(tmp_icb_cmd_ready_130), 
    .i_dat(tmp_icb_cmd_pack_130),
    .o_vld(tmp_icb_cmd_valid_131), 
    .o_rdy(delay_stage_select[131] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_131), 
    .o_dat(tmp_icb_cmd_pack_131),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_132;
  wire     tmp_icb_cmd_valid_132;
  wire     tmp_icb_cmd_ready_132;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_132 (
    .i_vld(tmp_icb_cmd_valid_131), 
    .i_rdy(tmp_icb_cmd_ready_131), 
    .i_dat(tmp_icb_cmd_pack_131),
    .o_vld(tmp_icb_cmd_valid_132), 
    .o_rdy(delay_stage_select[132] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_132), 
    .o_dat(tmp_icb_cmd_pack_132),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_133;
  wire     tmp_icb_cmd_valid_133;
  wire     tmp_icb_cmd_ready_133;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_133 (
    .i_vld(tmp_icb_cmd_valid_132), 
    .i_rdy(tmp_icb_cmd_ready_132), 
    .i_dat(tmp_icb_cmd_pack_132),
    .o_vld(tmp_icb_cmd_valid_133), 
    .o_rdy(delay_stage_select[133] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_133), 
    .o_dat(tmp_icb_cmd_pack_133),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_134;
  wire     tmp_icb_cmd_valid_134;
  wire     tmp_icb_cmd_ready_134;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_134 (
    .i_vld(tmp_icb_cmd_valid_133), 
    .i_rdy(tmp_icb_cmd_ready_133), 
    .i_dat(tmp_icb_cmd_pack_133),
    .o_vld(tmp_icb_cmd_valid_134), 
    .o_rdy(delay_stage_select[134] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_134), 
    .o_dat(tmp_icb_cmd_pack_134),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_135;
  wire     tmp_icb_cmd_valid_135;
  wire     tmp_icb_cmd_ready_135;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_135 (
    .i_vld(tmp_icb_cmd_valid_134), 
    .i_rdy(tmp_icb_cmd_ready_134), 
    .i_dat(tmp_icb_cmd_pack_134),
    .o_vld(tmp_icb_cmd_valid_135), 
    .o_rdy(delay_stage_select[135] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_135), 
    .o_dat(tmp_icb_cmd_pack_135),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_136;
  wire     tmp_icb_cmd_valid_136;
  wire     tmp_icb_cmd_ready_136;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_136 (
    .i_vld(tmp_icb_cmd_valid_135), 
    .i_rdy(tmp_icb_cmd_ready_135), 
    .i_dat(tmp_icb_cmd_pack_135),
    .o_vld(tmp_icb_cmd_valid_136), 
    .o_rdy(delay_stage_select[136] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_136), 
    .o_dat(tmp_icb_cmd_pack_136),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_137;
  wire     tmp_icb_cmd_valid_137;
  wire     tmp_icb_cmd_ready_137;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_137 (
    .i_vld(tmp_icb_cmd_valid_136), 
    .i_rdy(tmp_icb_cmd_ready_136), 
    .i_dat(tmp_icb_cmd_pack_136),
    .o_vld(tmp_icb_cmd_valid_137), 
    .o_rdy(delay_stage_select[137] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_137), 
    .o_dat(tmp_icb_cmd_pack_137),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_138;
  wire     tmp_icb_cmd_valid_138;
  wire     tmp_icb_cmd_ready_138;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_138 (
    .i_vld(tmp_icb_cmd_valid_137), 
    .i_rdy(tmp_icb_cmd_ready_137), 
    .i_dat(tmp_icb_cmd_pack_137),
    .o_vld(tmp_icb_cmd_valid_138), 
    .o_rdy(delay_stage_select[138] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_138), 
    .o_dat(tmp_icb_cmd_pack_138),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_139;
  wire     tmp_icb_cmd_valid_139;
  wire     tmp_icb_cmd_ready_139;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_139 (
    .i_vld(tmp_icb_cmd_valid_138), 
    .i_rdy(tmp_icb_cmd_ready_138), 
    .i_dat(tmp_icb_cmd_pack_138),
    .o_vld(tmp_icb_cmd_valid_139), 
    .o_rdy(delay_stage_select[139] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_139), 
    .o_dat(tmp_icb_cmd_pack_139),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_140;
  wire     tmp_icb_cmd_valid_140;
  wire     tmp_icb_cmd_ready_140;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_140 (
    .i_vld(tmp_icb_cmd_valid_139), 
    .i_rdy(tmp_icb_cmd_ready_139), 
    .i_dat(tmp_icb_cmd_pack_139),
    .o_vld(tmp_icb_cmd_valid_140), 
    .o_rdy(delay_stage_select[140] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_140), 
    .o_dat(tmp_icb_cmd_pack_140),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_141;
  wire     tmp_icb_cmd_valid_141;
  wire     tmp_icb_cmd_ready_141;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_141 (
    .i_vld(tmp_icb_cmd_valid_140), 
    .i_rdy(tmp_icb_cmd_ready_140), 
    .i_dat(tmp_icb_cmd_pack_140),
    .o_vld(tmp_icb_cmd_valid_141), 
    .o_rdy(delay_stage_select[141] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_141), 
    .o_dat(tmp_icb_cmd_pack_141),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_142;
  wire     tmp_icb_cmd_valid_142;
  wire     tmp_icb_cmd_ready_142;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_142 (
    .i_vld(tmp_icb_cmd_valid_141), 
    .i_rdy(tmp_icb_cmd_ready_141), 
    .i_dat(tmp_icb_cmd_pack_141),
    .o_vld(tmp_icb_cmd_valid_142), 
    .o_rdy(delay_stage_select[142] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_142), 
    .o_dat(tmp_icb_cmd_pack_142),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_143;
  wire     tmp_icb_cmd_valid_143;
  wire     tmp_icb_cmd_ready_143;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_143 (
    .i_vld(tmp_icb_cmd_valid_142), 
    .i_rdy(tmp_icb_cmd_ready_142), 
    .i_dat(tmp_icb_cmd_pack_142),
    .o_vld(tmp_icb_cmd_valid_143), 
    .o_rdy(delay_stage_select[143] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_143), 
    .o_dat(tmp_icb_cmd_pack_143),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_144;
  wire     tmp_icb_cmd_valid_144;
  wire     tmp_icb_cmd_ready_144;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_144 (
    .i_vld(tmp_icb_cmd_valid_143), 
    .i_rdy(tmp_icb_cmd_ready_143), 
    .i_dat(tmp_icb_cmd_pack_143),
    .o_vld(tmp_icb_cmd_valid_144), 
    .o_rdy(delay_stage_select[144] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_144), 
    .o_dat(tmp_icb_cmd_pack_144),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_145;
  wire     tmp_icb_cmd_valid_145;
  wire     tmp_icb_cmd_ready_145;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_145 (
    .i_vld(tmp_icb_cmd_valid_144), 
    .i_rdy(tmp_icb_cmd_ready_144), 
    .i_dat(tmp_icb_cmd_pack_144),
    .o_vld(tmp_icb_cmd_valid_145), 
    .o_rdy(delay_stage_select[145] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_145), 
    .o_dat(tmp_icb_cmd_pack_145),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_146;
  wire     tmp_icb_cmd_valid_146;
  wire     tmp_icb_cmd_ready_146;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_146 (
    .i_vld(tmp_icb_cmd_valid_145), 
    .i_rdy(tmp_icb_cmd_ready_145), 
    .i_dat(tmp_icb_cmd_pack_145),
    .o_vld(tmp_icb_cmd_valid_146), 
    .o_rdy(delay_stage_select[146] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_146), 
    .o_dat(tmp_icb_cmd_pack_146),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_147;
  wire     tmp_icb_cmd_valid_147;
  wire     tmp_icb_cmd_ready_147;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_147 (
    .i_vld(tmp_icb_cmd_valid_146), 
    .i_rdy(tmp_icb_cmd_ready_146), 
    .i_dat(tmp_icb_cmd_pack_146),
    .o_vld(tmp_icb_cmd_valid_147), 
    .o_rdy(delay_stage_select[147] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_147), 
    .o_dat(tmp_icb_cmd_pack_147),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_148;
  wire     tmp_icb_cmd_valid_148;
  wire     tmp_icb_cmd_ready_148;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_148 (
    .i_vld(tmp_icb_cmd_valid_147), 
    .i_rdy(tmp_icb_cmd_ready_147), 
    .i_dat(tmp_icb_cmd_pack_147),
    .o_vld(tmp_icb_cmd_valid_148), 
    .o_rdy(delay_stage_select[148] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_148), 
    .o_dat(tmp_icb_cmd_pack_148),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_149;
  wire     tmp_icb_cmd_valid_149;
  wire     tmp_icb_cmd_ready_149;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_149 (
    .i_vld(tmp_icb_cmd_valid_148), 
    .i_rdy(tmp_icb_cmd_ready_148), 
    .i_dat(tmp_icb_cmd_pack_148),
    .o_vld(tmp_icb_cmd_valid_149), 
    .o_rdy(delay_stage_select[149] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_149), 
    .o_dat(tmp_icb_cmd_pack_149),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_150;
  wire     tmp_icb_cmd_valid_150;
  wire     tmp_icb_cmd_ready_150;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_150 (
    .i_vld(tmp_icb_cmd_valid_149), 
    .i_rdy(tmp_icb_cmd_ready_149), 
    .i_dat(tmp_icb_cmd_pack_149),
    .o_vld(tmp_icb_cmd_valid_150), 
    .o_rdy(delay_stage_select[150] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_150), 
    .o_dat(tmp_icb_cmd_pack_150),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_151;
  wire     tmp_icb_cmd_valid_151;
  wire     tmp_icb_cmd_ready_151;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_151 (
    .i_vld(tmp_icb_cmd_valid_150), 
    .i_rdy(tmp_icb_cmd_ready_150), 
    .i_dat(tmp_icb_cmd_pack_150),
    .o_vld(tmp_icb_cmd_valid_151), 
    .o_rdy(delay_stage_select[151] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_151), 
    .o_dat(tmp_icb_cmd_pack_151),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_152;
  wire     tmp_icb_cmd_valid_152;
  wire     tmp_icb_cmd_ready_152;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_152 (
    .i_vld(tmp_icb_cmd_valid_151), 
    .i_rdy(tmp_icb_cmd_ready_151), 
    .i_dat(tmp_icb_cmd_pack_151),
    .o_vld(tmp_icb_cmd_valid_152), 
    .o_rdy(delay_stage_select[152] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_152), 
    .o_dat(tmp_icb_cmd_pack_152),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_153;
  wire     tmp_icb_cmd_valid_153;
  wire     tmp_icb_cmd_ready_153;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_153 (
    .i_vld(tmp_icb_cmd_valid_152), 
    .i_rdy(tmp_icb_cmd_ready_152), 
    .i_dat(tmp_icb_cmd_pack_152),
    .o_vld(tmp_icb_cmd_valid_153), 
    .o_rdy(delay_stage_select[153] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_153), 
    .o_dat(tmp_icb_cmd_pack_153),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_154;
  wire     tmp_icb_cmd_valid_154;
  wire     tmp_icb_cmd_ready_154;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_154 (
    .i_vld(tmp_icb_cmd_valid_153), 
    .i_rdy(tmp_icb_cmd_ready_153), 
    .i_dat(tmp_icb_cmd_pack_153),
    .o_vld(tmp_icb_cmd_valid_154), 
    .o_rdy(delay_stage_select[154] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_154), 
    .o_dat(tmp_icb_cmd_pack_154),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_155;
  wire     tmp_icb_cmd_valid_155;
  wire     tmp_icb_cmd_ready_155;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_155 (
    .i_vld(tmp_icb_cmd_valid_154), 
    .i_rdy(tmp_icb_cmd_ready_154), 
    .i_dat(tmp_icb_cmd_pack_154),
    .o_vld(tmp_icb_cmd_valid_155), 
    .o_rdy(delay_stage_select[155] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_155), 
    .o_dat(tmp_icb_cmd_pack_155),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_156;
  wire     tmp_icb_cmd_valid_156;
  wire     tmp_icb_cmd_ready_156;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_156 (
    .i_vld(tmp_icb_cmd_valid_155), 
    .i_rdy(tmp_icb_cmd_ready_155), 
    .i_dat(tmp_icb_cmd_pack_155),
    .o_vld(tmp_icb_cmd_valid_156), 
    .o_rdy(delay_stage_select[156] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_156), 
    .o_dat(tmp_icb_cmd_pack_156),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_157;
  wire     tmp_icb_cmd_valid_157;
  wire     tmp_icb_cmd_ready_157;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_157 (
    .i_vld(tmp_icb_cmd_valid_156), 
    .i_rdy(tmp_icb_cmd_ready_156), 
    .i_dat(tmp_icb_cmd_pack_156),
    .o_vld(tmp_icb_cmd_valid_157), 
    .o_rdy(delay_stage_select[157] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_157), 
    .o_dat(tmp_icb_cmd_pack_157),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_158;
  wire     tmp_icb_cmd_valid_158;
  wire     tmp_icb_cmd_ready_158;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_158 (
    .i_vld(tmp_icb_cmd_valid_157), 
    .i_rdy(tmp_icb_cmd_ready_157), 
    .i_dat(tmp_icb_cmd_pack_157),
    .o_vld(tmp_icb_cmd_valid_158), 
    .o_rdy(delay_stage_select[158] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_158), 
    .o_dat(tmp_icb_cmd_pack_158),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_159;
  wire     tmp_icb_cmd_valid_159;
  wire     tmp_icb_cmd_ready_159;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_159 (
    .i_vld(tmp_icb_cmd_valid_158), 
    .i_rdy(tmp_icb_cmd_ready_158), 
    .i_dat(tmp_icb_cmd_pack_158),
    .o_vld(tmp_icb_cmd_valid_159), 
    .o_rdy(delay_stage_select[159] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_159), 
    .o_dat(tmp_icb_cmd_pack_159),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_160;
  wire     tmp_icb_cmd_valid_160;
  wire     tmp_icb_cmd_ready_160;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_160 (
    .i_vld(tmp_icb_cmd_valid_159), 
    .i_rdy(tmp_icb_cmd_ready_159), 
    .i_dat(tmp_icb_cmd_pack_159),
    .o_vld(tmp_icb_cmd_valid_160), 
    .o_rdy(delay_stage_select[160] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_160), 
    .o_dat(tmp_icb_cmd_pack_160),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_161;
  wire     tmp_icb_cmd_valid_161;
  wire     tmp_icb_cmd_ready_161;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_161 (
    .i_vld(tmp_icb_cmd_valid_160), 
    .i_rdy(tmp_icb_cmd_ready_160), 
    .i_dat(tmp_icb_cmd_pack_160),
    .o_vld(tmp_icb_cmd_valid_161), 
    .o_rdy(delay_stage_select[161] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_161), 
    .o_dat(tmp_icb_cmd_pack_161),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_162;
  wire     tmp_icb_cmd_valid_162;
  wire     tmp_icb_cmd_ready_162;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_162 (
    .i_vld(tmp_icb_cmd_valid_161), 
    .i_rdy(tmp_icb_cmd_ready_161), 
    .i_dat(tmp_icb_cmd_pack_161),
    .o_vld(tmp_icb_cmd_valid_162), 
    .o_rdy(delay_stage_select[162] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_162), 
    .o_dat(tmp_icb_cmd_pack_162),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_163;
  wire     tmp_icb_cmd_valid_163;
  wire     tmp_icb_cmd_ready_163;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_163 (
    .i_vld(tmp_icb_cmd_valid_162), 
    .i_rdy(tmp_icb_cmd_ready_162), 
    .i_dat(tmp_icb_cmd_pack_162),
    .o_vld(tmp_icb_cmd_valid_163), 
    .o_rdy(delay_stage_select[163] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_163), 
    .o_dat(tmp_icb_cmd_pack_163),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_164;
  wire     tmp_icb_cmd_valid_164;
  wire     tmp_icb_cmd_ready_164;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_164 (
    .i_vld(tmp_icb_cmd_valid_163), 
    .i_rdy(tmp_icb_cmd_ready_163), 
    .i_dat(tmp_icb_cmd_pack_163),
    .o_vld(tmp_icb_cmd_valid_164), 
    .o_rdy(delay_stage_select[164] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_164), 
    .o_dat(tmp_icb_cmd_pack_164),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_165;
  wire     tmp_icb_cmd_valid_165;
  wire     tmp_icb_cmd_ready_165;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_165 (
    .i_vld(tmp_icb_cmd_valid_164), 
    .i_rdy(tmp_icb_cmd_ready_164), 
    .i_dat(tmp_icb_cmd_pack_164),
    .o_vld(tmp_icb_cmd_valid_165), 
    .o_rdy(delay_stage_select[165] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_165), 
    .o_dat(tmp_icb_cmd_pack_165),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_166;
  wire     tmp_icb_cmd_valid_166;
  wire     tmp_icb_cmd_ready_166;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_166 (
    .i_vld(tmp_icb_cmd_valid_165), 
    .i_rdy(tmp_icb_cmd_ready_165), 
    .i_dat(tmp_icb_cmd_pack_165),
    .o_vld(tmp_icb_cmd_valid_166), 
    .o_rdy(delay_stage_select[166] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_166), 
    .o_dat(tmp_icb_cmd_pack_166),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_167;
  wire     tmp_icb_cmd_valid_167;
  wire     tmp_icb_cmd_ready_167;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_167 (
    .i_vld(tmp_icb_cmd_valid_166), 
    .i_rdy(tmp_icb_cmd_ready_166), 
    .i_dat(tmp_icb_cmd_pack_166),
    .o_vld(tmp_icb_cmd_valid_167), 
    .o_rdy(delay_stage_select[167] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_167), 
    .o_dat(tmp_icb_cmd_pack_167),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_168;
  wire     tmp_icb_cmd_valid_168;
  wire     tmp_icb_cmd_ready_168;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_168 (
    .i_vld(tmp_icb_cmd_valid_167), 
    .i_rdy(tmp_icb_cmd_ready_167), 
    .i_dat(tmp_icb_cmd_pack_167),
    .o_vld(tmp_icb_cmd_valid_168), 
    .o_rdy(delay_stage_select[168] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_168), 
    .o_dat(tmp_icb_cmd_pack_168),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_169;
  wire     tmp_icb_cmd_valid_169;
  wire     tmp_icb_cmd_ready_169;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_169 (
    .i_vld(tmp_icb_cmd_valid_168), 
    .i_rdy(tmp_icb_cmd_ready_168), 
    .i_dat(tmp_icb_cmd_pack_168),
    .o_vld(tmp_icb_cmd_valid_169), 
    .o_rdy(delay_stage_select[169] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_169), 
    .o_dat(tmp_icb_cmd_pack_169),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_170;
  wire     tmp_icb_cmd_valid_170;
  wire     tmp_icb_cmd_ready_170;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_170 (
    .i_vld(tmp_icb_cmd_valid_169), 
    .i_rdy(tmp_icb_cmd_ready_169), 
    .i_dat(tmp_icb_cmd_pack_169),
    .o_vld(tmp_icb_cmd_valid_170), 
    .o_rdy(delay_stage_select[170] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_170), 
    .o_dat(tmp_icb_cmd_pack_170),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_171;
  wire     tmp_icb_cmd_valid_171;
  wire     tmp_icb_cmd_ready_171;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_171 (
    .i_vld(tmp_icb_cmd_valid_170), 
    .i_rdy(tmp_icb_cmd_ready_170), 
    .i_dat(tmp_icb_cmd_pack_170),
    .o_vld(tmp_icb_cmd_valid_171), 
    .o_rdy(delay_stage_select[171] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_171), 
    .o_dat(tmp_icb_cmd_pack_171),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_172;
  wire     tmp_icb_cmd_valid_172;
  wire     tmp_icb_cmd_ready_172;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_172 (
    .i_vld(tmp_icb_cmd_valid_171), 
    .i_rdy(tmp_icb_cmd_ready_171), 
    .i_dat(tmp_icb_cmd_pack_171),
    .o_vld(tmp_icb_cmd_valid_172), 
    .o_rdy(delay_stage_select[172] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_172), 
    .o_dat(tmp_icb_cmd_pack_172),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_173;
  wire     tmp_icb_cmd_valid_173;
  wire     tmp_icb_cmd_ready_173;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_173 (
    .i_vld(tmp_icb_cmd_valid_172), 
    .i_rdy(tmp_icb_cmd_ready_172), 
    .i_dat(tmp_icb_cmd_pack_172),
    .o_vld(tmp_icb_cmd_valid_173), 
    .o_rdy(delay_stage_select[173] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_173), 
    .o_dat(tmp_icb_cmd_pack_173),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_174;
  wire     tmp_icb_cmd_valid_174;
  wire     tmp_icb_cmd_ready_174;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_174 (
    .i_vld(tmp_icb_cmd_valid_173), 
    .i_rdy(tmp_icb_cmd_ready_173), 
    .i_dat(tmp_icb_cmd_pack_173),
    .o_vld(tmp_icb_cmd_valid_174), 
    .o_rdy(delay_stage_select[174] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_174), 
    .o_dat(tmp_icb_cmd_pack_174),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_175;
  wire     tmp_icb_cmd_valid_175;
  wire     tmp_icb_cmd_ready_175;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_175 (
    .i_vld(tmp_icb_cmd_valid_174), 
    .i_rdy(tmp_icb_cmd_ready_174), 
    .i_dat(tmp_icb_cmd_pack_174),
    .o_vld(tmp_icb_cmd_valid_175), 
    .o_rdy(delay_stage_select[175] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_175), 
    .o_dat(tmp_icb_cmd_pack_175),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_176;
  wire     tmp_icb_cmd_valid_176;
  wire     tmp_icb_cmd_ready_176;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_176 (
    .i_vld(tmp_icb_cmd_valid_175), 
    .i_rdy(tmp_icb_cmd_ready_175), 
    .i_dat(tmp_icb_cmd_pack_175),
    .o_vld(tmp_icb_cmd_valid_176), 
    .o_rdy(delay_stage_select[176] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_176), 
    .o_dat(tmp_icb_cmd_pack_176),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_177;
  wire     tmp_icb_cmd_valid_177;
  wire     tmp_icb_cmd_ready_177;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_177 (
    .i_vld(tmp_icb_cmd_valid_176), 
    .i_rdy(tmp_icb_cmd_ready_176), 
    .i_dat(tmp_icb_cmd_pack_176),
    .o_vld(tmp_icb_cmd_valid_177), 
    .o_rdy(delay_stage_select[177] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_177), 
    .o_dat(tmp_icb_cmd_pack_177),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_178;
  wire     tmp_icb_cmd_valid_178;
  wire     tmp_icb_cmd_ready_178;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_178 (
    .i_vld(tmp_icb_cmd_valid_177), 
    .i_rdy(tmp_icb_cmd_ready_177), 
    .i_dat(tmp_icb_cmd_pack_177),
    .o_vld(tmp_icb_cmd_valid_178), 
    .o_rdy(delay_stage_select[178] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_178), 
    .o_dat(tmp_icb_cmd_pack_178),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_179;
  wire     tmp_icb_cmd_valid_179;
  wire     tmp_icb_cmd_ready_179;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_179 (
    .i_vld(tmp_icb_cmd_valid_178), 
    .i_rdy(tmp_icb_cmd_ready_178), 
    .i_dat(tmp_icb_cmd_pack_178),
    .o_vld(tmp_icb_cmd_valid_179), 
    .o_rdy(delay_stage_select[179] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_179), 
    .o_dat(tmp_icb_cmd_pack_179),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_180;
  wire     tmp_icb_cmd_valid_180;
  wire     tmp_icb_cmd_ready_180;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_180 (
    .i_vld(tmp_icb_cmd_valid_179), 
    .i_rdy(tmp_icb_cmd_ready_179), 
    .i_dat(tmp_icb_cmd_pack_179),
    .o_vld(tmp_icb_cmd_valid_180), 
    .o_rdy(delay_stage_select[180] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_180), 
    .o_dat(tmp_icb_cmd_pack_180),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_181;
  wire     tmp_icb_cmd_valid_181;
  wire     tmp_icb_cmd_ready_181;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_181 (
    .i_vld(tmp_icb_cmd_valid_180), 
    .i_rdy(tmp_icb_cmd_ready_180), 
    .i_dat(tmp_icb_cmd_pack_180),
    .o_vld(tmp_icb_cmd_valid_181), 
    .o_rdy(delay_stage_select[181] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_181), 
    .o_dat(tmp_icb_cmd_pack_181),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_182;
  wire     tmp_icb_cmd_valid_182;
  wire     tmp_icb_cmd_ready_182;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_182 (
    .i_vld(tmp_icb_cmd_valid_181), 
    .i_rdy(tmp_icb_cmd_ready_181), 
    .i_dat(tmp_icb_cmd_pack_181),
    .o_vld(tmp_icb_cmd_valid_182), 
    .o_rdy(delay_stage_select[182] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_182), 
    .o_dat(tmp_icb_cmd_pack_182),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_183;
  wire     tmp_icb_cmd_valid_183;
  wire     tmp_icb_cmd_ready_183;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_183 (
    .i_vld(tmp_icb_cmd_valid_182), 
    .i_rdy(tmp_icb_cmd_ready_182), 
    .i_dat(tmp_icb_cmd_pack_182),
    .o_vld(tmp_icb_cmd_valid_183), 
    .o_rdy(delay_stage_select[183] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_183), 
    .o_dat(tmp_icb_cmd_pack_183),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_184;
  wire     tmp_icb_cmd_valid_184;
  wire     tmp_icb_cmd_ready_184;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_184 (
    .i_vld(tmp_icb_cmd_valid_183), 
    .i_rdy(tmp_icb_cmd_ready_183), 
    .i_dat(tmp_icb_cmd_pack_183),
    .o_vld(tmp_icb_cmd_valid_184), 
    .o_rdy(delay_stage_select[184] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_184), 
    .o_dat(tmp_icb_cmd_pack_184),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_185;
  wire     tmp_icb_cmd_valid_185;
  wire     tmp_icb_cmd_ready_185;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_185 (
    .i_vld(tmp_icb_cmd_valid_184), 
    .i_rdy(tmp_icb_cmd_ready_184), 
    .i_dat(tmp_icb_cmd_pack_184),
    .o_vld(tmp_icb_cmd_valid_185), 
    .o_rdy(delay_stage_select[185] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_185), 
    .o_dat(tmp_icb_cmd_pack_185),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_186;
  wire     tmp_icb_cmd_valid_186;
  wire     tmp_icb_cmd_ready_186;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_186 (
    .i_vld(tmp_icb_cmd_valid_185), 
    .i_rdy(tmp_icb_cmd_ready_185), 
    .i_dat(tmp_icb_cmd_pack_185),
    .o_vld(tmp_icb_cmd_valid_186), 
    .o_rdy(delay_stage_select[186] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_186), 
    .o_dat(tmp_icb_cmd_pack_186),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_187;
  wire     tmp_icb_cmd_valid_187;
  wire     tmp_icb_cmd_ready_187;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_187 (
    .i_vld(tmp_icb_cmd_valid_186), 
    .i_rdy(tmp_icb_cmd_ready_186), 
    .i_dat(tmp_icb_cmd_pack_186),
    .o_vld(tmp_icb_cmd_valid_187), 
    .o_rdy(delay_stage_select[187] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_187), 
    .o_dat(tmp_icb_cmd_pack_187),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_188;
  wire     tmp_icb_cmd_valid_188;
  wire     tmp_icb_cmd_ready_188;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_188 (
    .i_vld(tmp_icb_cmd_valid_187), 
    .i_rdy(tmp_icb_cmd_ready_187), 
    .i_dat(tmp_icb_cmd_pack_187),
    .o_vld(tmp_icb_cmd_valid_188), 
    .o_rdy(delay_stage_select[188] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_188), 
    .o_dat(tmp_icb_cmd_pack_188),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_189;
  wire     tmp_icb_cmd_valid_189;
  wire     tmp_icb_cmd_ready_189;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_189 (
    .i_vld(tmp_icb_cmd_valid_188), 
    .i_rdy(tmp_icb_cmd_ready_188), 
    .i_dat(tmp_icb_cmd_pack_188),
    .o_vld(tmp_icb_cmd_valid_189), 
    .o_rdy(delay_stage_select[189] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_189), 
    .o_dat(tmp_icb_cmd_pack_189),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_190;
  wire     tmp_icb_cmd_valid_190;
  wire     tmp_icb_cmd_ready_190;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_190 (
    .i_vld(tmp_icb_cmd_valid_189), 
    .i_rdy(tmp_icb_cmd_ready_189), 
    .i_dat(tmp_icb_cmd_pack_189),
    .o_vld(tmp_icb_cmd_valid_190), 
    .o_rdy(delay_stage_select[190] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_190), 
    .o_dat(tmp_icb_cmd_pack_190),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_191;
  wire     tmp_icb_cmd_valid_191;
  wire     tmp_icb_cmd_ready_191;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_191 (
    .i_vld(tmp_icb_cmd_valid_190), 
    .i_rdy(tmp_icb_cmd_ready_190), 
    .i_dat(tmp_icb_cmd_pack_190),
    .o_vld(tmp_icb_cmd_valid_191), 
    .o_rdy(delay_stage_select[191] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_191), 
    .o_dat(tmp_icb_cmd_pack_191),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_192;
  wire     tmp_icb_cmd_valid_192;
  wire     tmp_icb_cmd_ready_192;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_192 (
    .i_vld(tmp_icb_cmd_valid_191), 
    .i_rdy(tmp_icb_cmd_ready_191), 
    .i_dat(tmp_icb_cmd_pack_191),
    .o_vld(tmp_icb_cmd_valid_192), 
    .o_rdy(delay_stage_select[192] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_192), 
    .o_dat(tmp_icb_cmd_pack_192),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_193;
  wire     tmp_icb_cmd_valid_193;
  wire     tmp_icb_cmd_ready_193;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_193 (
    .i_vld(tmp_icb_cmd_valid_192), 
    .i_rdy(tmp_icb_cmd_ready_192), 
    .i_dat(tmp_icb_cmd_pack_192),
    .o_vld(tmp_icb_cmd_valid_193), 
    .o_rdy(delay_stage_select[193] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_193), 
    .o_dat(tmp_icb_cmd_pack_193),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_194;
  wire     tmp_icb_cmd_valid_194;
  wire     tmp_icb_cmd_ready_194;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_194 (
    .i_vld(tmp_icb_cmd_valid_193), 
    .i_rdy(tmp_icb_cmd_ready_193), 
    .i_dat(tmp_icb_cmd_pack_193),
    .o_vld(tmp_icb_cmd_valid_194), 
    .o_rdy(delay_stage_select[194] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_194), 
    .o_dat(tmp_icb_cmd_pack_194),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_195;
  wire     tmp_icb_cmd_valid_195;
  wire     tmp_icb_cmd_ready_195;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_195 (
    .i_vld(tmp_icb_cmd_valid_194), 
    .i_rdy(tmp_icb_cmd_ready_194), 
    .i_dat(tmp_icb_cmd_pack_194),
    .o_vld(tmp_icb_cmd_valid_195), 
    .o_rdy(delay_stage_select[195] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_195), 
    .o_dat(tmp_icb_cmd_pack_195),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_196;
  wire     tmp_icb_cmd_valid_196;
  wire     tmp_icb_cmd_ready_196;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_196 (
    .i_vld(tmp_icb_cmd_valid_195), 
    .i_rdy(tmp_icb_cmd_ready_195), 
    .i_dat(tmp_icb_cmd_pack_195),
    .o_vld(tmp_icb_cmd_valid_196), 
    .o_rdy(delay_stage_select[196] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_196), 
    .o_dat(tmp_icb_cmd_pack_196),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_197;
  wire     tmp_icb_cmd_valid_197;
  wire     tmp_icb_cmd_ready_197;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_197 (
    .i_vld(tmp_icb_cmd_valid_196), 
    .i_rdy(tmp_icb_cmd_ready_196), 
    .i_dat(tmp_icb_cmd_pack_196),
    .o_vld(tmp_icb_cmd_valid_197), 
    .o_rdy(delay_stage_select[197] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_197), 
    .o_dat(tmp_icb_cmd_pack_197),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_198;
  wire     tmp_icb_cmd_valid_198;
  wire     tmp_icb_cmd_ready_198;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_198 (
    .i_vld(tmp_icb_cmd_valid_197), 
    .i_rdy(tmp_icb_cmd_ready_197), 
    .i_dat(tmp_icb_cmd_pack_197),
    .o_vld(tmp_icb_cmd_valid_198), 
    .o_rdy(delay_stage_select[198] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_198), 
    .o_dat(tmp_icb_cmd_pack_198),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_199;
  wire     tmp_icb_cmd_valid_199;
  wire     tmp_icb_cmd_ready_199;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_199 (
    .i_vld(tmp_icb_cmd_valid_198), 
    .i_rdy(tmp_icb_cmd_ready_198), 
    .i_dat(tmp_icb_cmd_pack_198),
    .o_vld(tmp_icb_cmd_valid_199), 
    .o_rdy(delay_stage_select[199] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_199), 
    .o_dat(tmp_icb_cmd_pack_199),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_200;
  wire     tmp_icb_cmd_valid_200;
  wire     tmp_icb_cmd_ready_200;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_200 (
    .i_vld(tmp_icb_cmd_valid_199), 
    .i_rdy(tmp_icb_cmd_ready_199), 
    .i_dat(tmp_icb_cmd_pack_199),
    .o_vld(tmp_icb_cmd_valid_200), 
    .o_rdy(delay_stage_select[200] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_200), 
    .o_dat(tmp_icb_cmd_pack_200),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_201;
  wire     tmp_icb_cmd_valid_201;
  wire     tmp_icb_cmd_ready_201;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_201 (
    .i_vld(tmp_icb_cmd_valid_200), 
    .i_rdy(tmp_icb_cmd_ready_200), 
    .i_dat(tmp_icb_cmd_pack_200),
    .o_vld(tmp_icb_cmd_valid_201), 
    .o_rdy(delay_stage_select[201] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_201), 
    .o_dat(tmp_icb_cmd_pack_201),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_202;
  wire     tmp_icb_cmd_valid_202;
  wire     tmp_icb_cmd_ready_202;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_202 (
    .i_vld(tmp_icb_cmd_valid_201), 
    .i_rdy(tmp_icb_cmd_ready_201), 
    .i_dat(tmp_icb_cmd_pack_201),
    .o_vld(tmp_icb_cmd_valid_202), 
    .o_rdy(delay_stage_select[202] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_202), 
    .o_dat(tmp_icb_cmd_pack_202),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_203;
  wire     tmp_icb_cmd_valid_203;
  wire     tmp_icb_cmd_ready_203;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_203 (
    .i_vld(tmp_icb_cmd_valid_202), 
    .i_rdy(tmp_icb_cmd_ready_202), 
    .i_dat(tmp_icb_cmd_pack_202),
    .o_vld(tmp_icb_cmd_valid_203), 
    .o_rdy(delay_stage_select[203] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_203), 
    .o_dat(tmp_icb_cmd_pack_203),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_204;
  wire     tmp_icb_cmd_valid_204;
  wire     tmp_icb_cmd_ready_204;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_204 (
    .i_vld(tmp_icb_cmd_valid_203), 
    .i_rdy(tmp_icb_cmd_ready_203), 
    .i_dat(tmp_icb_cmd_pack_203),
    .o_vld(tmp_icb_cmd_valid_204), 
    .o_rdy(delay_stage_select[204] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_204), 
    .o_dat(tmp_icb_cmd_pack_204),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_205;
  wire     tmp_icb_cmd_valid_205;
  wire     tmp_icb_cmd_ready_205;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_205 (
    .i_vld(tmp_icb_cmd_valid_204), 
    .i_rdy(tmp_icb_cmd_ready_204), 
    .i_dat(tmp_icb_cmd_pack_204),
    .o_vld(tmp_icb_cmd_valid_205), 
    .o_rdy(delay_stage_select[205] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_205), 
    .o_dat(tmp_icb_cmd_pack_205),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_206;
  wire     tmp_icb_cmd_valid_206;
  wire     tmp_icb_cmd_ready_206;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_206 (
    .i_vld(tmp_icb_cmd_valid_205), 
    .i_rdy(tmp_icb_cmd_ready_205), 
    .i_dat(tmp_icb_cmd_pack_205),
    .o_vld(tmp_icb_cmd_valid_206), 
    .o_rdy(delay_stage_select[206] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_206), 
    .o_dat(tmp_icb_cmd_pack_206),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_207;
  wire     tmp_icb_cmd_valid_207;
  wire     tmp_icb_cmd_ready_207;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_207 (
    .i_vld(tmp_icb_cmd_valid_206), 
    .i_rdy(tmp_icb_cmd_ready_206), 
    .i_dat(tmp_icb_cmd_pack_206),
    .o_vld(tmp_icb_cmd_valid_207), 
    .o_rdy(delay_stage_select[207] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_207), 
    .o_dat(tmp_icb_cmd_pack_207),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_208;
  wire     tmp_icb_cmd_valid_208;
  wire     tmp_icb_cmd_ready_208;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_208 (
    .i_vld(tmp_icb_cmd_valid_207), 
    .i_rdy(tmp_icb_cmd_ready_207), 
    .i_dat(tmp_icb_cmd_pack_207),
    .o_vld(tmp_icb_cmd_valid_208), 
    .o_rdy(delay_stage_select[208] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_208), 
    .o_dat(tmp_icb_cmd_pack_208),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_209;
  wire     tmp_icb_cmd_valid_209;
  wire     tmp_icb_cmd_ready_209;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_209 (
    .i_vld(tmp_icb_cmd_valid_208), 
    .i_rdy(tmp_icb_cmd_ready_208), 
    .i_dat(tmp_icb_cmd_pack_208),
    .o_vld(tmp_icb_cmd_valid_209), 
    .o_rdy(delay_stage_select[209] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_209), 
    .o_dat(tmp_icb_cmd_pack_209),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_210;
  wire     tmp_icb_cmd_valid_210;
  wire     tmp_icb_cmd_ready_210;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_210 (
    .i_vld(tmp_icb_cmd_valid_209), 
    .i_rdy(tmp_icb_cmd_ready_209), 
    .i_dat(tmp_icb_cmd_pack_209),
    .o_vld(tmp_icb_cmd_valid_210), 
    .o_rdy(delay_stage_select[210] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_210), 
    .o_dat(tmp_icb_cmd_pack_210),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_211;
  wire     tmp_icb_cmd_valid_211;
  wire     tmp_icb_cmd_ready_211;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_211 (
    .i_vld(tmp_icb_cmd_valid_210), 
    .i_rdy(tmp_icb_cmd_ready_210), 
    .i_dat(tmp_icb_cmd_pack_210),
    .o_vld(tmp_icb_cmd_valid_211), 
    .o_rdy(delay_stage_select[211] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_211), 
    .o_dat(tmp_icb_cmd_pack_211),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_212;
  wire     tmp_icb_cmd_valid_212;
  wire     tmp_icb_cmd_ready_212;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_212 (
    .i_vld(tmp_icb_cmd_valid_211), 
    .i_rdy(tmp_icb_cmd_ready_211), 
    .i_dat(tmp_icb_cmd_pack_211),
    .o_vld(tmp_icb_cmd_valid_212), 
    .o_rdy(delay_stage_select[212] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_212), 
    .o_dat(tmp_icb_cmd_pack_212),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_213;
  wire     tmp_icb_cmd_valid_213;
  wire     tmp_icb_cmd_ready_213;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_213 (
    .i_vld(tmp_icb_cmd_valid_212), 
    .i_rdy(tmp_icb_cmd_ready_212), 
    .i_dat(tmp_icb_cmd_pack_212),
    .o_vld(tmp_icb_cmd_valid_213), 
    .o_rdy(delay_stage_select[213] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_213), 
    .o_dat(tmp_icb_cmd_pack_213),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_214;
  wire     tmp_icb_cmd_valid_214;
  wire     tmp_icb_cmd_ready_214;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_214 (
    .i_vld(tmp_icb_cmd_valid_213), 
    .i_rdy(tmp_icb_cmd_ready_213), 
    .i_dat(tmp_icb_cmd_pack_213),
    .o_vld(tmp_icb_cmd_valid_214), 
    .o_rdy(delay_stage_select[214] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_214), 
    .o_dat(tmp_icb_cmd_pack_214),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_215;
  wire     tmp_icb_cmd_valid_215;
  wire     tmp_icb_cmd_ready_215;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_215 (
    .i_vld(tmp_icb_cmd_valid_214), 
    .i_rdy(tmp_icb_cmd_ready_214), 
    .i_dat(tmp_icb_cmd_pack_214),
    .o_vld(tmp_icb_cmd_valid_215), 
    .o_rdy(delay_stage_select[215] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_215), 
    .o_dat(tmp_icb_cmd_pack_215),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_216;
  wire     tmp_icb_cmd_valid_216;
  wire     tmp_icb_cmd_ready_216;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_216 (
    .i_vld(tmp_icb_cmd_valid_215), 
    .i_rdy(tmp_icb_cmd_ready_215), 
    .i_dat(tmp_icb_cmd_pack_215),
    .o_vld(tmp_icb_cmd_valid_216), 
    .o_rdy(delay_stage_select[216] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_216), 
    .o_dat(tmp_icb_cmd_pack_216),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_217;
  wire     tmp_icb_cmd_valid_217;
  wire     tmp_icb_cmd_ready_217;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_217 (
    .i_vld(tmp_icb_cmd_valid_216), 
    .i_rdy(tmp_icb_cmd_ready_216), 
    .i_dat(tmp_icb_cmd_pack_216),
    .o_vld(tmp_icb_cmd_valid_217), 
    .o_rdy(delay_stage_select[217] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_217), 
    .o_dat(tmp_icb_cmd_pack_217),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_218;
  wire     tmp_icb_cmd_valid_218;
  wire     tmp_icb_cmd_ready_218;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_218 (
    .i_vld(tmp_icb_cmd_valid_217), 
    .i_rdy(tmp_icb_cmd_ready_217), 
    .i_dat(tmp_icb_cmd_pack_217),
    .o_vld(tmp_icb_cmd_valid_218), 
    .o_rdy(delay_stage_select[218] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_218), 
    .o_dat(tmp_icb_cmd_pack_218),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_219;
  wire     tmp_icb_cmd_valid_219;
  wire     tmp_icb_cmd_ready_219;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_219 (
    .i_vld(tmp_icb_cmd_valid_218), 
    .i_rdy(tmp_icb_cmd_ready_218), 
    .i_dat(tmp_icb_cmd_pack_218),
    .o_vld(tmp_icb_cmd_valid_219), 
    .o_rdy(delay_stage_select[219] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_219), 
    .o_dat(tmp_icb_cmd_pack_219),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_220;
  wire     tmp_icb_cmd_valid_220;
  wire     tmp_icb_cmd_ready_220;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_220 (
    .i_vld(tmp_icb_cmd_valid_219), 
    .i_rdy(tmp_icb_cmd_ready_219), 
    .i_dat(tmp_icb_cmd_pack_219),
    .o_vld(tmp_icb_cmd_valid_220), 
    .o_rdy(delay_stage_select[220] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_220), 
    .o_dat(tmp_icb_cmd_pack_220),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_221;
  wire     tmp_icb_cmd_valid_221;
  wire     tmp_icb_cmd_ready_221;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_221 (
    .i_vld(tmp_icb_cmd_valid_220), 
    .i_rdy(tmp_icb_cmd_ready_220), 
    .i_dat(tmp_icb_cmd_pack_220),
    .o_vld(tmp_icb_cmd_valid_221), 
    .o_rdy(delay_stage_select[221] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_221), 
    .o_dat(tmp_icb_cmd_pack_221),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_222;
  wire     tmp_icb_cmd_valid_222;
  wire     tmp_icb_cmd_ready_222;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_222 (
    .i_vld(tmp_icb_cmd_valid_221), 
    .i_rdy(tmp_icb_cmd_ready_221), 
    .i_dat(tmp_icb_cmd_pack_221),
    .o_vld(tmp_icb_cmd_valid_222), 
    .o_rdy(delay_stage_select[222] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_222), 
    .o_dat(tmp_icb_cmd_pack_222),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_223;
  wire     tmp_icb_cmd_valid_223;
  wire     tmp_icb_cmd_ready_223;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_223 (
    .i_vld(tmp_icb_cmd_valid_222), 
    .i_rdy(tmp_icb_cmd_ready_222), 
    .i_dat(tmp_icb_cmd_pack_222),
    .o_vld(tmp_icb_cmd_valid_223), 
    .o_rdy(delay_stage_select[223] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_223), 
    .o_dat(tmp_icb_cmd_pack_223),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_224;
  wire     tmp_icb_cmd_valid_224;
  wire     tmp_icb_cmd_ready_224;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_224 (
    .i_vld(tmp_icb_cmd_valid_223), 
    .i_rdy(tmp_icb_cmd_ready_223), 
    .i_dat(tmp_icb_cmd_pack_223),
    .o_vld(tmp_icb_cmd_valid_224), 
    .o_rdy(delay_stage_select[224] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_224), 
    .o_dat(tmp_icb_cmd_pack_224),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_225;
  wire     tmp_icb_cmd_valid_225;
  wire     tmp_icb_cmd_ready_225;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_225 (
    .i_vld(tmp_icb_cmd_valid_224), 
    .i_rdy(tmp_icb_cmd_ready_224), 
    .i_dat(tmp_icb_cmd_pack_224),
    .o_vld(tmp_icb_cmd_valid_225), 
    .o_rdy(delay_stage_select[225] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_225), 
    .o_dat(tmp_icb_cmd_pack_225),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_226;
  wire     tmp_icb_cmd_valid_226;
  wire     tmp_icb_cmd_ready_226;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_226 (
    .i_vld(tmp_icb_cmd_valid_225), 
    .i_rdy(tmp_icb_cmd_ready_225), 
    .i_dat(tmp_icb_cmd_pack_225),
    .o_vld(tmp_icb_cmd_valid_226), 
    .o_rdy(delay_stage_select[226] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_226), 
    .o_dat(tmp_icb_cmd_pack_226),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_227;
  wire     tmp_icb_cmd_valid_227;
  wire     tmp_icb_cmd_ready_227;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_227 (
    .i_vld(tmp_icb_cmd_valid_226), 
    .i_rdy(tmp_icb_cmd_ready_226), 
    .i_dat(tmp_icb_cmd_pack_226),
    .o_vld(tmp_icb_cmd_valid_227), 
    .o_rdy(delay_stage_select[227] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_227), 
    .o_dat(tmp_icb_cmd_pack_227),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_228;
  wire     tmp_icb_cmd_valid_228;
  wire     tmp_icb_cmd_ready_228;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_228 (
    .i_vld(tmp_icb_cmd_valid_227), 
    .i_rdy(tmp_icb_cmd_ready_227), 
    .i_dat(tmp_icb_cmd_pack_227),
    .o_vld(tmp_icb_cmd_valid_228), 
    .o_rdy(delay_stage_select[228] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_228), 
    .o_dat(tmp_icb_cmd_pack_228),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_229;
  wire     tmp_icb_cmd_valid_229;
  wire     tmp_icb_cmd_ready_229;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_229 (
    .i_vld(tmp_icb_cmd_valid_228), 
    .i_rdy(tmp_icb_cmd_ready_228), 
    .i_dat(tmp_icb_cmd_pack_228),
    .o_vld(tmp_icb_cmd_valid_229), 
    .o_rdy(delay_stage_select[229] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_229), 
    .o_dat(tmp_icb_cmd_pack_229),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_230;
  wire     tmp_icb_cmd_valid_230;
  wire     tmp_icb_cmd_ready_230;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_230 (
    .i_vld(tmp_icb_cmd_valid_229), 
    .i_rdy(tmp_icb_cmd_ready_229), 
    .i_dat(tmp_icb_cmd_pack_229),
    .o_vld(tmp_icb_cmd_valid_230), 
    .o_rdy(delay_stage_select[230] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_230), 
    .o_dat(tmp_icb_cmd_pack_230),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_231;
  wire     tmp_icb_cmd_valid_231;
  wire     tmp_icb_cmd_ready_231;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_231 (
    .i_vld(tmp_icb_cmd_valid_230), 
    .i_rdy(tmp_icb_cmd_ready_230), 
    .i_dat(tmp_icb_cmd_pack_230),
    .o_vld(tmp_icb_cmd_valid_231), 
    .o_rdy(delay_stage_select[231] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_231), 
    .o_dat(tmp_icb_cmd_pack_231),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_232;
  wire     tmp_icb_cmd_valid_232;
  wire     tmp_icb_cmd_ready_232;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_232 (
    .i_vld(tmp_icb_cmd_valid_231), 
    .i_rdy(tmp_icb_cmd_ready_231), 
    .i_dat(tmp_icb_cmd_pack_231),
    .o_vld(tmp_icb_cmd_valid_232), 
    .o_rdy(delay_stage_select[232] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_232), 
    .o_dat(tmp_icb_cmd_pack_232),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_233;
  wire     tmp_icb_cmd_valid_233;
  wire     tmp_icb_cmd_ready_233;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_233 (
    .i_vld(tmp_icb_cmd_valid_232), 
    .i_rdy(tmp_icb_cmd_ready_232), 
    .i_dat(tmp_icb_cmd_pack_232),
    .o_vld(tmp_icb_cmd_valid_233), 
    .o_rdy(delay_stage_select[233] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_233), 
    .o_dat(tmp_icb_cmd_pack_233),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_234;
  wire     tmp_icb_cmd_valid_234;
  wire     tmp_icb_cmd_ready_234;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_234 (
    .i_vld(tmp_icb_cmd_valid_233), 
    .i_rdy(tmp_icb_cmd_ready_233), 
    .i_dat(tmp_icb_cmd_pack_233),
    .o_vld(tmp_icb_cmd_valid_234), 
    .o_rdy(delay_stage_select[234] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_234), 
    .o_dat(tmp_icb_cmd_pack_234),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_235;
  wire     tmp_icb_cmd_valid_235;
  wire     tmp_icb_cmd_ready_235;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_235 (
    .i_vld(tmp_icb_cmd_valid_234), 
    .i_rdy(tmp_icb_cmd_ready_234), 
    .i_dat(tmp_icb_cmd_pack_234),
    .o_vld(tmp_icb_cmd_valid_235), 
    .o_rdy(delay_stage_select[235] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_235), 
    .o_dat(tmp_icb_cmd_pack_235),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_236;
  wire     tmp_icb_cmd_valid_236;
  wire     tmp_icb_cmd_ready_236;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_236 (
    .i_vld(tmp_icb_cmd_valid_235), 
    .i_rdy(tmp_icb_cmd_ready_235), 
    .i_dat(tmp_icb_cmd_pack_235),
    .o_vld(tmp_icb_cmd_valid_236), 
    .o_rdy(delay_stage_select[236] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_236), 
    .o_dat(tmp_icb_cmd_pack_236),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_237;
  wire     tmp_icb_cmd_valid_237;
  wire     tmp_icb_cmd_ready_237;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_237 (
    .i_vld(tmp_icb_cmd_valid_236), 
    .i_rdy(tmp_icb_cmd_ready_236), 
    .i_dat(tmp_icb_cmd_pack_236),
    .o_vld(tmp_icb_cmd_valid_237), 
    .o_rdy(delay_stage_select[237] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_237), 
    .o_dat(tmp_icb_cmd_pack_237),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_238;
  wire     tmp_icb_cmd_valid_238;
  wire     tmp_icb_cmd_ready_238;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_238 (
    .i_vld(tmp_icb_cmd_valid_237), 
    .i_rdy(tmp_icb_cmd_ready_237), 
    .i_dat(tmp_icb_cmd_pack_237),
    .o_vld(tmp_icb_cmd_valid_238), 
    .o_rdy(delay_stage_select[238] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_238), 
    .o_dat(tmp_icb_cmd_pack_238),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_239;
  wire     tmp_icb_cmd_valid_239;
  wire     tmp_icb_cmd_ready_239;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_239 (
    .i_vld(tmp_icb_cmd_valid_238), 
    .i_rdy(tmp_icb_cmd_ready_238), 
    .i_dat(tmp_icb_cmd_pack_238),
    .o_vld(tmp_icb_cmd_valid_239), 
    .o_rdy(delay_stage_select[239] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_239), 
    .o_dat(tmp_icb_cmd_pack_239),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_240;
  wire     tmp_icb_cmd_valid_240;
  wire     tmp_icb_cmd_ready_240;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_240 (
    .i_vld(tmp_icb_cmd_valid_239), 
    .i_rdy(tmp_icb_cmd_ready_239), 
    .i_dat(tmp_icb_cmd_pack_239),
    .o_vld(tmp_icb_cmd_valid_240), 
    .o_rdy(delay_stage_select[240] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_240), 
    .o_dat(tmp_icb_cmd_pack_240),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_241;
  wire     tmp_icb_cmd_valid_241;
  wire     tmp_icb_cmd_ready_241;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_241 (
    .i_vld(tmp_icb_cmd_valid_240), 
    .i_rdy(tmp_icb_cmd_ready_240), 
    .i_dat(tmp_icb_cmd_pack_240),
    .o_vld(tmp_icb_cmd_valid_241), 
    .o_rdy(delay_stage_select[241] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_241), 
    .o_dat(tmp_icb_cmd_pack_241),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_242;
  wire     tmp_icb_cmd_valid_242;
  wire     tmp_icb_cmd_ready_242;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_242 (
    .i_vld(tmp_icb_cmd_valid_241), 
    .i_rdy(tmp_icb_cmd_ready_241), 
    .i_dat(tmp_icb_cmd_pack_241),
    .o_vld(tmp_icb_cmd_valid_242), 
    .o_rdy(delay_stage_select[242] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_242), 
    .o_dat(tmp_icb_cmd_pack_242),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_243;
  wire     tmp_icb_cmd_valid_243;
  wire     tmp_icb_cmd_ready_243;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_243 (
    .i_vld(tmp_icb_cmd_valid_242), 
    .i_rdy(tmp_icb_cmd_ready_242), 
    .i_dat(tmp_icb_cmd_pack_242),
    .o_vld(tmp_icb_cmd_valid_243), 
    .o_rdy(delay_stage_select[243] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_243), 
    .o_dat(tmp_icb_cmd_pack_243),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_244;
  wire     tmp_icb_cmd_valid_244;
  wire     tmp_icb_cmd_ready_244;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_244 (
    .i_vld(tmp_icb_cmd_valid_243), 
    .i_rdy(tmp_icb_cmd_ready_243), 
    .i_dat(tmp_icb_cmd_pack_243),
    .o_vld(tmp_icb_cmd_valid_244), 
    .o_rdy(delay_stage_select[244] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_244), 
    .o_dat(tmp_icb_cmd_pack_244),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_245;
  wire     tmp_icb_cmd_valid_245;
  wire     tmp_icb_cmd_ready_245;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_245 (
    .i_vld(tmp_icb_cmd_valid_244), 
    .i_rdy(tmp_icb_cmd_ready_244), 
    .i_dat(tmp_icb_cmd_pack_244),
    .o_vld(tmp_icb_cmd_valid_245), 
    .o_rdy(delay_stage_select[245] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_245), 
    .o_dat(tmp_icb_cmd_pack_245),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_246;
  wire     tmp_icb_cmd_valid_246;
  wire     tmp_icb_cmd_ready_246;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_246 (
    .i_vld(tmp_icb_cmd_valid_245), 
    .i_rdy(tmp_icb_cmd_ready_245), 
    .i_dat(tmp_icb_cmd_pack_245),
    .o_vld(tmp_icb_cmd_valid_246), 
    .o_rdy(delay_stage_select[246] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_246), 
    .o_dat(tmp_icb_cmd_pack_246),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_247;
  wire     tmp_icb_cmd_valid_247;
  wire     tmp_icb_cmd_ready_247;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_247 (
    .i_vld(tmp_icb_cmd_valid_246), 
    .i_rdy(tmp_icb_cmd_ready_246), 
    .i_dat(tmp_icb_cmd_pack_246),
    .o_vld(tmp_icb_cmd_valid_247), 
    .o_rdy(delay_stage_select[247] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_247), 
    .o_dat(tmp_icb_cmd_pack_247),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_248;
  wire     tmp_icb_cmd_valid_248;
  wire     tmp_icb_cmd_ready_248;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_248 (
    .i_vld(tmp_icb_cmd_valid_247), 
    .i_rdy(tmp_icb_cmd_ready_247), 
    .i_dat(tmp_icb_cmd_pack_247),
    .o_vld(tmp_icb_cmd_valid_248), 
    .o_rdy(delay_stage_select[248] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_248), 
    .o_dat(tmp_icb_cmd_pack_248),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_249;
  wire     tmp_icb_cmd_valid_249;
  wire     tmp_icb_cmd_ready_249;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_249 (
    .i_vld(tmp_icb_cmd_valid_248), 
    .i_rdy(tmp_icb_cmd_ready_248), 
    .i_dat(tmp_icb_cmd_pack_248),
    .o_vld(tmp_icb_cmd_valid_249), 
    .o_rdy(delay_stage_select[249] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_249), 
    .o_dat(tmp_icb_cmd_pack_249),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_250;
  wire     tmp_icb_cmd_valid_250;
  wire     tmp_icb_cmd_ready_250;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_250 (
    .i_vld(tmp_icb_cmd_valid_249), 
    .i_rdy(tmp_icb_cmd_ready_249), 
    .i_dat(tmp_icb_cmd_pack_249),
    .o_vld(tmp_icb_cmd_valid_250), 
    .o_rdy(delay_stage_select[250] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_250), 
    .o_dat(tmp_icb_cmd_pack_250),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_251;
  wire     tmp_icb_cmd_valid_251;
  wire     tmp_icb_cmd_ready_251;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_251 (
    .i_vld(tmp_icb_cmd_valid_250), 
    .i_rdy(tmp_icb_cmd_ready_250), 
    .i_dat(tmp_icb_cmd_pack_250),
    .o_vld(tmp_icb_cmd_valid_251), 
    .o_rdy(delay_stage_select[251] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_251), 
    .o_dat(tmp_icb_cmd_pack_251),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_252;
  wire     tmp_icb_cmd_valid_252;
  wire     tmp_icb_cmd_ready_252;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_252 (
    .i_vld(tmp_icb_cmd_valid_251), 
    .i_rdy(tmp_icb_cmd_ready_251), 
    .i_dat(tmp_icb_cmd_pack_251),
    .o_vld(tmp_icb_cmd_valid_252), 
    .o_rdy(delay_stage_select[252] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_252), 
    .o_dat(tmp_icb_cmd_pack_252),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_253;
  wire     tmp_icb_cmd_valid_253;
  wire     tmp_icb_cmd_ready_253;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_253 (
    .i_vld(tmp_icb_cmd_valid_252), 
    .i_rdy(tmp_icb_cmd_ready_252), 
    .i_dat(tmp_icb_cmd_pack_252),
    .o_vld(tmp_icb_cmd_valid_253), 
    .o_rdy(delay_stage_select[253] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_253), 
    .o_dat(tmp_icb_cmd_pack_253),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_254;
  wire     tmp_icb_cmd_valid_254;
  wire     tmp_icb_cmd_ready_254;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_254 (
    .i_vld(tmp_icb_cmd_valid_253), 
    .i_rdy(tmp_icb_cmd_ready_253), 
    .i_dat(tmp_icb_cmd_pack_253),
    .o_vld(tmp_icb_cmd_valid_254), 
    .o_rdy(delay_stage_select[254] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_254), 
    .o_dat(tmp_icb_cmd_pack_254),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_255;
  wire     tmp_icb_cmd_valid_255;
  wire     tmp_icb_cmd_ready_255;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_255 (
    .i_vld(tmp_icb_cmd_valid_254), 
    .i_rdy(tmp_icb_cmd_ready_254), 
    .i_dat(tmp_icb_cmd_pack_254),
    .o_vld(tmp_icb_cmd_valid_255), 
    .o_rdy(delay_stage_select[255] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_255), 
    .o_dat(tmp_icb_cmd_pack_255),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_256;
  wire     tmp_icb_cmd_valid_256;
  wire     tmp_icb_cmd_ready_256;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_256 (
    .i_vld(tmp_icb_cmd_valid_255), 
    .i_rdy(tmp_icb_cmd_ready_255), 
    .i_dat(tmp_icb_cmd_pack_255),
    .o_vld(tmp_icb_cmd_valid_256), 
    .o_rdy(delay_stage_select[256] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_256), 
    .o_dat(tmp_icb_cmd_pack_256),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_257;
  wire     tmp_icb_cmd_valid_257;
  wire     tmp_icb_cmd_ready_257;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_257 (
    .i_vld(tmp_icb_cmd_valid_256), 
    .i_rdy(tmp_icb_cmd_ready_256), 
    .i_dat(tmp_icb_cmd_pack_256),
    .o_vld(tmp_icb_cmd_valid_257), 
    .o_rdy(delay_stage_select[257] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_257), 
    .o_dat(tmp_icb_cmd_pack_257),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_258;
  wire     tmp_icb_cmd_valid_258;
  wire     tmp_icb_cmd_ready_258;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_258 (
    .i_vld(tmp_icb_cmd_valid_257), 
    .i_rdy(tmp_icb_cmd_ready_257), 
    .i_dat(tmp_icb_cmd_pack_257),
    .o_vld(tmp_icb_cmd_valid_258), 
    .o_rdy(delay_stage_select[258] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_258), 
    .o_dat(tmp_icb_cmd_pack_258),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_259;
  wire     tmp_icb_cmd_valid_259;
  wire     tmp_icb_cmd_ready_259;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_259 (
    .i_vld(tmp_icb_cmd_valid_258), 
    .i_rdy(tmp_icb_cmd_ready_258), 
    .i_dat(tmp_icb_cmd_pack_258),
    .o_vld(tmp_icb_cmd_valid_259), 
    .o_rdy(delay_stage_select[259] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_259), 
    .o_dat(tmp_icb_cmd_pack_259),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_260;
  wire     tmp_icb_cmd_valid_260;
  wire     tmp_icb_cmd_ready_260;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_260 (
    .i_vld(tmp_icb_cmd_valid_259), 
    .i_rdy(tmp_icb_cmd_ready_259), 
    .i_dat(tmp_icb_cmd_pack_259),
    .o_vld(tmp_icb_cmd_valid_260), 
    .o_rdy(delay_stage_select[260] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_260), 
    .o_dat(tmp_icb_cmd_pack_260),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_261;
  wire     tmp_icb_cmd_valid_261;
  wire     tmp_icb_cmd_ready_261;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_261 (
    .i_vld(tmp_icb_cmd_valid_260), 
    .i_rdy(tmp_icb_cmd_ready_260), 
    .i_dat(tmp_icb_cmd_pack_260),
    .o_vld(tmp_icb_cmd_valid_261), 
    .o_rdy(delay_stage_select[261] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_261), 
    .o_dat(tmp_icb_cmd_pack_261),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_262;
  wire     tmp_icb_cmd_valid_262;
  wire     tmp_icb_cmd_ready_262;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_262 (
    .i_vld(tmp_icb_cmd_valid_261), 
    .i_rdy(tmp_icb_cmd_ready_261), 
    .i_dat(tmp_icb_cmd_pack_261),
    .o_vld(tmp_icb_cmd_valid_262), 
    .o_rdy(delay_stage_select[262] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_262), 
    .o_dat(tmp_icb_cmd_pack_262),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_263;
  wire     tmp_icb_cmd_valid_263;
  wire     tmp_icb_cmd_ready_263;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_263 (
    .i_vld(tmp_icb_cmd_valid_262), 
    .i_rdy(tmp_icb_cmd_ready_262), 
    .i_dat(tmp_icb_cmd_pack_262),
    .o_vld(tmp_icb_cmd_valid_263), 
    .o_rdy(delay_stage_select[263] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_263), 
    .o_dat(tmp_icb_cmd_pack_263),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_264;
  wire     tmp_icb_cmd_valid_264;
  wire     tmp_icb_cmd_ready_264;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_264 (
    .i_vld(tmp_icb_cmd_valid_263), 
    .i_rdy(tmp_icb_cmd_ready_263), 
    .i_dat(tmp_icb_cmd_pack_263),
    .o_vld(tmp_icb_cmd_valid_264), 
    .o_rdy(delay_stage_select[264] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_264), 
    .o_dat(tmp_icb_cmd_pack_264),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_265;
  wire     tmp_icb_cmd_valid_265;
  wire     tmp_icb_cmd_ready_265;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_265 (
    .i_vld(tmp_icb_cmd_valid_264), 
    .i_rdy(tmp_icb_cmd_ready_264), 
    .i_dat(tmp_icb_cmd_pack_264),
    .o_vld(tmp_icb_cmd_valid_265), 
    .o_rdy(delay_stage_select[265] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_265), 
    .o_dat(tmp_icb_cmd_pack_265),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_266;
  wire     tmp_icb_cmd_valid_266;
  wire     tmp_icb_cmd_ready_266;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_266 (
    .i_vld(tmp_icb_cmd_valid_265), 
    .i_rdy(tmp_icb_cmd_ready_265), 
    .i_dat(tmp_icb_cmd_pack_265),
    .o_vld(tmp_icb_cmd_valid_266), 
    .o_rdy(delay_stage_select[266] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_266), 
    .o_dat(tmp_icb_cmd_pack_266),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_267;
  wire     tmp_icb_cmd_valid_267;
  wire     tmp_icb_cmd_ready_267;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_267 (
    .i_vld(tmp_icb_cmd_valid_266), 
    .i_rdy(tmp_icb_cmd_ready_266), 
    .i_dat(tmp_icb_cmd_pack_266),
    .o_vld(tmp_icb_cmd_valid_267), 
    .o_rdy(delay_stage_select[267] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_267), 
    .o_dat(tmp_icb_cmd_pack_267),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_268;
  wire     tmp_icb_cmd_valid_268;
  wire     tmp_icb_cmd_ready_268;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_268 (
    .i_vld(tmp_icb_cmd_valid_267), 
    .i_rdy(tmp_icb_cmd_ready_267), 
    .i_dat(tmp_icb_cmd_pack_267),
    .o_vld(tmp_icb_cmd_valid_268), 
    .o_rdy(delay_stage_select[268] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_268), 
    .o_dat(tmp_icb_cmd_pack_268),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_269;
  wire     tmp_icb_cmd_valid_269;
  wire     tmp_icb_cmd_ready_269;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_269 (
    .i_vld(tmp_icb_cmd_valid_268), 
    .i_rdy(tmp_icb_cmd_ready_268), 
    .i_dat(tmp_icb_cmd_pack_268),
    .o_vld(tmp_icb_cmd_valid_269), 
    .o_rdy(delay_stage_select[269] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_269), 
    .o_dat(tmp_icb_cmd_pack_269),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_270;
  wire     tmp_icb_cmd_valid_270;
  wire     tmp_icb_cmd_ready_270;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_270 (
    .i_vld(tmp_icb_cmd_valid_269), 
    .i_rdy(tmp_icb_cmd_ready_269), 
    .i_dat(tmp_icb_cmd_pack_269),
    .o_vld(tmp_icb_cmd_valid_270), 
    .o_rdy(delay_stage_select[270] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_270), 
    .o_dat(tmp_icb_cmd_pack_270),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_271;
  wire     tmp_icb_cmd_valid_271;
  wire     tmp_icb_cmd_ready_271;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_271 (
    .i_vld(tmp_icb_cmd_valid_270), 
    .i_rdy(tmp_icb_cmd_ready_270), 
    .i_dat(tmp_icb_cmd_pack_270),
    .o_vld(tmp_icb_cmd_valid_271), 
    .o_rdy(delay_stage_select[271] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_271), 
    .o_dat(tmp_icb_cmd_pack_271),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_272;
  wire     tmp_icb_cmd_valid_272;
  wire     tmp_icb_cmd_ready_272;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_272 (
    .i_vld(tmp_icb_cmd_valid_271), 
    .i_rdy(tmp_icb_cmd_ready_271), 
    .i_dat(tmp_icb_cmd_pack_271),
    .o_vld(tmp_icb_cmd_valid_272), 
    .o_rdy(delay_stage_select[272] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_272), 
    .o_dat(tmp_icb_cmd_pack_272),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_273;
  wire     tmp_icb_cmd_valid_273;
  wire     tmp_icb_cmd_ready_273;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_273 (
    .i_vld(tmp_icb_cmd_valid_272), 
    .i_rdy(tmp_icb_cmd_ready_272), 
    .i_dat(tmp_icb_cmd_pack_272),
    .o_vld(tmp_icb_cmd_valid_273), 
    .o_rdy(delay_stage_select[273] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_273), 
    .o_dat(tmp_icb_cmd_pack_273),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_274;
  wire     tmp_icb_cmd_valid_274;
  wire     tmp_icb_cmd_ready_274;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_274 (
    .i_vld(tmp_icb_cmd_valid_273), 
    .i_rdy(tmp_icb_cmd_ready_273), 
    .i_dat(tmp_icb_cmd_pack_273),
    .o_vld(tmp_icb_cmd_valid_274), 
    .o_rdy(delay_stage_select[274] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_274), 
    .o_dat(tmp_icb_cmd_pack_274),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_275;
  wire     tmp_icb_cmd_valid_275;
  wire     tmp_icb_cmd_ready_275;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_275 (
    .i_vld(tmp_icb_cmd_valid_274), 
    .i_rdy(tmp_icb_cmd_ready_274), 
    .i_dat(tmp_icb_cmd_pack_274),
    .o_vld(tmp_icb_cmd_valid_275), 
    .o_rdy(delay_stage_select[275] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_275), 
    .o_dat(tmp_icb_cmd_pack_275),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_276;
  wire     tmp_icb_cmd_valid_276;
  wire     tmp_icb_cmd_ready_276;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_276 (
    .i_vld(tmp_icb_cmd_valid_275), 
    .i_rdy(tmp_icb_cmd_ready_275), 
    .i_dat(tmp_icb_cmd_pack_275),
    .o_vld(tmp_icb_cmd_valid_276), 
    .o_rdy(delay_stage_select[276] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_276), 
    .o_dat(tmp_icb_cmd_pack_276),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_277;
  wire     tmp_icb_cmd_valid_277;
  wire     tmp_icb_cmd_ready_277;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_277 (
    .i_vld(tmp_icb_cmd_valid_276), 
    .i_rdy(tmp_icb_cmd_ready_276), 
    .i_dat(tmp_icb_cmd_pack_276),
    .o_vld(tmp_icb_cmd_valid_277), 
    .o_rdy(delay_stage_select[277] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_277), 
    .o_dat(tmp_icb_cmd_pack_277),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_278;
  wire     tmp_icb_cmd_valid_278;
  wire     tmp_icb_cmd_ready_278;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_278 (
    .i_vld(tmp_icb_cmd_valid_277), 
    .i_rdy(tmp_icb_cmd_ready_277), 
    .i_dat(tmp_icb_cmd_pack_277),
    .o_vld(tmp_icb_cmd_valid_278), 
    .o_rdy(delay_stage_select[278] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_278), 
    .o_dat(tmp_icb_cmd_pack_278),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_279;
  wire     tmp_icb_cmd_valid_279;
  wire     tmp_icb_cmd_ready_279;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_279 (
    .i_vld(tmp_icb_cmd_valid_278), 
    .i_rdy(tmp_icb_cmd_ready_278), 
    .i_dat(tmp_icb_cmd_pack_278),
    .o_vld(tmp_icb_cmd_valid_279), 
    .o_rdy(delay_stage_select[279] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_279), 
    .o_dat(tmp_icb_cmd_pack_279),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_280;
  wire     tmp_icb_cmd_valid_280;
  wire     tmp_icb_cmd_ready_280;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_280 (
    .i_vld(tmp_icb_cmd_valid_279), 
    .i_rdy(tmp_icb_cmd_ready_279), 
    .i_dat(tmp_icb_cmd_pack_279),
    .o_vld(tmp_icb_cmd_valid_280), 
    .o_rdy(delay_stage_select[280] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_280), 
    .o_dat(tmp_icb_cmd_pack_280),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_281;
  wire     tmp_icb_cmd_valid_281;
  wire     tmp_icb_cmd_ready_281;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_281 (
    .i_vld(tmp_icb_cmd_valid_280), 
    .i_rdy(tmp_icb_cmd_ready_280), 
    .i_dat(tmp_icb_cmd_pack_280),
    .o_vld(tmp_icb_cmd_valid_281), 
    .o_rdy(delay_stage_select[281] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_281), 
    .o_dat(tmp_icb_cmd_pack_281),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_282;
  wire     tmp_icb_cmd_valid_282;
  wire     tmp_icb_cmd_ready_282;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_282 (
    .i_vld(tmp_icb_cmd_valid_281), 
    .i_rdy(tmp_icb_cmd_ready_281), 
    .i_dat(tmp_icb_cmd_pack_281),
    .o_vld(tmp_icb_cmd_valid_282), 
    .o_rdy(delay_stage_select[282] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_282), 
    .o_dat(tmp_icb_cmd_pack_282),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_283;
  wire     tmp_icb_cmd_valid_283;
  wire     tmp_icb_cmd_ready_283;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_283 (
    .i_vld(tmp_icb_cmd_valid_282), 
    .i_rdy(tmp_icb_cmd_ready_282), 
    .i_dat(tmp_icb_cmd_pack_282),
    .o_vld(tmp_icb_cmd_valid_283), 
    .o_rdy(delay_stage_select[283] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_283), 
    .o_dat(tmp_icb_cmd_pack_283),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_284;
  wire     tmp_icb_cmd_valid_284;
  wire     tmp_icb_cmd_ready_284;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_284 (
    .i_vld(tmp_icb_cmd_valid_283), 
    .i_rdy(tmp_icb_cmd_ready_283), 
    .i_dat(tmp_icb_cmd_pack_283),
    .o_vld(tmp_icb_cmd_valid_284), 
    .o_rdy(delay_stage_select[284] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_284), 
    .o_dat(tmp_icb_cmd_pack_284),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_285;
  wire     tmp_icb_cmd_valid_285;
  wire     tmp_icb_cmd_ready_285;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_285 (
    .i_vld(tmp_icb_cmd_valid_284), 
    .i_rdy(tmp_icb_cmd_ready_284), 
    .i_dat(tmp_icb_cmd_pack_284),
    .o_vld(tmp_icb_cmd_valid_285), 
    .o_rdy(delay_stage_select[285] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_285), 
    .o_dat(tmp_icb_cmd_pack_285),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_286;
  wire     tmp_icb_cmd_valid_286;
  wire     tmp_icb_cmd_ready_286;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_286 (
    .i_vld(tmp_icb_cmd_valid_285), 
    .i_rdy(tmp_icb_cmd_ready_285), 
    .i_dat(tmp_icb_cmd_pack_285),
    .o_vld(tmp_icb_cmd_valid_286), 
    .o_rdy(delay_stage_select[286] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_286), 
    .o_dat(tmp_icb_cmd_pack_286),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_287;
  wire     tmp_icb_cmd_valid_287;
  wire     tmp_icb_cmd_ready_287;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_287 (
    .i_vld(tmp_icb_cmd_valid_286), 
    .i_rdy(tmp_icb_cmd_ready_286), 
    .i_dat(tmp_icb_cmd_pack_286),
    .o_vld(tmp_icb_cmd_valid_287), 
    .o_rdy(delay_stage_select[287] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_287), 
    .o_dat(tmp_icb_cmd_pack_287),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_288;
  wire     tmp_icb_cmd_valid_288;
  wire     tmp_icb_cmd_ready_288;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_288 (
    .i_vld(tmp_icb_cmd_valid_287), 
    .i_rdy(tmp_icb_cmd_ready_287), 
    .i_dat(tmp_icb_cmd_pack_287),
    .o_vld(tmp_icb_cmd_valid_288), 
    .o_rdy(delay_stage_select[288] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_288), 
    .o_dat(tmp_icb_cmd_pack_288),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_289;
  wire     tmp_icb_cmd_valid_289;
  wire     tmp_icb_cmd_ready_289;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_289 (
    .i_vld(tmp_icb_cmd_valid_288), 
    .i_rdy(tmp_icb_cmd_ready_288), 
    .i_dat(tmp_icb_cmd_pack_288),
    .o_vld(tmp_icb_cmd_valid_289), 
    .o_rdy(delay_stage_select[289] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_289), 
    .o_dat(tmp_icb_cmd_pack_289),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_290;
  wire     tmp_icb_cmd_valid_290;
  wire     tmp_icb_cmd_ready_290;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_290 (
    .i_vld(tmp_icb_cmd_valid_289), 
    .i_rdy(tmp_icb_cmd_ready_289), 
    .i_dat(tmp_icb_cmd_pack_289),
    .o_vld(tmp_icb_cmd_valid_290), 
    .o_rdy(delay_stage_select[290] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_290), 
    .o_dat(tmp_icb_cmd_pack_290),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_291;
  wire     tmp_icb_cmd_valid_291;
  wire     tmp_icb_cmd_ready_291;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_291 (
    .i_vld(tmp_icb_cmd_valid_290), 
    .i_rdy(tmp_icb_cmd_ready_290), 
    .i_dat(tmp_icb_cmd_pack_290),
    .o_vld(tmp_icb_cmd_valid_291), 
    .o_rdy(delay_stage_select[291] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_291), 
    .o_dat(tmp_icb_cmd_pack_291),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_292;
  wire     tmp_icb_cmd_valid_292;
  wire     tmp_icb_cmd_ready_292;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_292 (
    .i_vld(tmp_icb_cmd_valid_291), 
    .i_rdy(tmp_icb_cmd_ready_291), 
    .i_dat(tmp_icb_cmd_pack_291),
    .o_vld(tmp_icb_cmd_valid_292), 
    .o_rdy(delay_stage_select[292] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_292), 
    .o_dat(tmp_icb_cmd_pack_292),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_293;
  wire     tmp_icb_cmd_valid_293;
  wire     tmp_icb_cmd_ready_293;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_293 (
    .i_vld(tmp_icb_cmd_valid_292), 
    .i_rdy(tmp_icb_cmd_ready_292), 
    .i_dat(tmp_icb_cmd_pack_292),
    .o_vld(tmp_icb_cmd_valid_293), 
    .o_rdy(delay_stage_select[293] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_293), 
    .o_dat(tmp_icb_cmd_pack_293),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_294;
  wire     tmp_icb_cmd_valid_294;
  wire     tmp_icb_cmd_ready_294;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_294 (
    .i_vld(tmp_icb_cmd_valid_293), 
    .i_rdy(tmp_icb_cmd_ready_293), 
    .i_dat(tmp_icb_cmd_pack_293),
    .o_vld(tmp_icb_cmd_valid_294), 
    .o_rdy(delay_stage_select[294] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_294), 
    .o_dat(tmp_icb_cmd_pack_294),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_295;
  wire     tmp_icb_cmd_valid_295;
  wire     tmp_icb_cmd_ready_295;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_295 (
    .i_vld(tmp_icb_cmd_valid_294), 
    .i_rdy(tmp_icb_cmd_ready_294), 
    .i_dat(tmp_icb_cmd_pack_294),
    .o_vld(tmp_icb_cmd_valid_295), 
    .o_rdy(delay_stage_select[295] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_295), 
    .o_dat(tmp_icb_cmd_pack_295),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_296;
  wire     tmp_icb_cmd_valid_296;
  wire     tmp_icb_cmd_ready_296;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_296 (
    .i_vld(tmp_icb_cmd_valid_295), 
    .i_rdy(tmp_icb_cmd_ready_295), 
    .i_dat(tmp_icb_cmd_pack_295),
    .o_vld(tmp_icb_cmd_valid_296), 
    .o_rdy(delay_stage_select[296] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_296), 
    .o_dat(tmp_icb_cmd_pack_296),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_297;
  wire     tmp_icb_cmd_valid_297;
  wire     tmp_icb_cmd_ready_297;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_297 (
    .i_vld(tmp_icb_cmd_valid_296), 
    .i_rdy(tmp_icb_cmd_ready_296), 
    .i_dat(tmp_icb_cmd_pack_296),
    .o_vld(tmp_icb_cmd_valid_297), 
    .o_rdy(delay_stage_select[297] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_297), 
    .o_dat(tmp_icb_cmd_pack_297),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_298;
  wire     tmp_icb_cmd_valid_298;
  wire     tmp_icb_cmd_ready_298;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_298 (
    .i_vld(tmp_icb_cmd_valid_297), 
    .i_rdy(tmp_icb_cmd_ready_297), 
    .i_dat(tmp_icb_cmd_pack_297),
    .o_vld(tmp_icb_cmd_valid_298), 
    .o_rdy(delay_stage_select[298] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_298), 
    .o_dat(tmp_icb_cmd_pack_298),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_299;
  wire     tmp_icb_cmd_valid_299;
  wire     tmp_icb_cmd_ready_299;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_299 (
    .i_vld(tmp_icb_cmd_valid_298), 
    .i_rdy(tmp_icb_cmd_ready_298), 
    .i_dat(tmp_icb_cmd_pack_298),
    .o_vld(tmp_icb_cmd_valid_299), 
    .o_rdy(delay_stage_select[299] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_299), 
    .o_dat(tmp_icb_cmd_pack_299),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_300;
  wire     tmp_icb_cmd_valid_300;
  wire     tmp_icb_cmd_ready_300;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_300 (
    .i_vld(tmp_icb_cmd_valid_299), 
    .i_rdy(tmp_icb_cmd_ready_299), 
    .i_dat(tmp_icb_cmd_pack_299),
    .o_vld(tmp_icb_cmd_valid_300), 
    .o_rdy(delay_stage_select[300] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_300), 
    .o_dat(tmp_icb_cmd_pack_300),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_301;
  wire     tmp_icb_cmd_valid_301;
  wire     tmp_icb_cmd_ready_301;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_301 (
    .i_vld(tmp_icb_cmd_valid_300), 
    .i_rdy(tmp_icb_cmd_ready_300), 
    .i_dat(tmp_icb_cmd_pack_300),
    .o_vld(tmp_icb_cmd_valid_301), 
    .o_rdy(delay_stage_select[301] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_301), 
    .o_dat(tmp_icb_cmd_pack_301),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_302;
  wire     tmp_icb_cmd_valid_302;
  wire     tmp_icb_cmd_ready_302;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_302 (
    .i_vld(tmp_icb_cmd_valid_301), 
    .i_rdy(tmp_icb_cmd_ready_301), 
    .i_dat(tmp_icb_cmd_pack_301),
    .o_vld(tmp_icb_cmd_valid_302), 
    .o_rdy(delay_stage_select[302] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_302), 
    .o_dat(tmp_icb_cmd_pack_302),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_303;
  wire     tmp_icb_cmd_valid_303;
  wire     tmp_icb_cmd_ready_303;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_303 (
    .i_vld(tmp_icb_cmd_valid_302), 
    .i_rdy(tmp_icb_cmd_ready_302), 
    .i_dat(tmp_icb_cmd_pack_302),
    .o_vld(tmp_icb_cmd_valid_303), 
    .o_rdy(delay_stage_select[303] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_303), 
    .o_dat(tmp_icb_cmd_pack_303),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_304;
  wire     tmp_icb_cmd_valid_304;
  wire     tmp_icb_cmd_ready_304;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_304 (
    .i_vld(tmp_icb_cmd_valid_303), 
    .i_rdy(tmp_icb_cmd_ready_303), 
    .i_dat(tmp_icb_cmd_pack_303),
    .o_vld(tmp_icb_cmd_valid_304), 
    .o_rdy(delay_stage_select[304] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_304), 
    .o_dat(tmp_icb_cmd_pack_304),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_305;
  wire     tmp_icb_cmd_valid_305;
  wire     tmp_icb_cmd_ready_305;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_305 (
    .i_vld(tmp_icb_cmd_valid_304), 
    .i_rdy(tmp_icb_cmd_ready_304), 
    .i_dat(tmp_icb_cmd_pack_304),
    .o_vld(tmp_icb_cmd_valid_305), 
    .o_rdy(delay_stage_select[305] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_305), 
    .o_dat(tmp_icb_cmd_pack_305),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_306;
  wire     tmp_icb_cmd_valid_306;
  wire     tmp_icb_cmd_ready_306;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_306 (
    .i_vld(tmp_icb_cmd_valid_305), 
    .i_rdy(tmp_icb_cmd_ready_305), 
    .i_dat(tmp_icb_cmd_pack_305),
    .o_vld(tmp_icb_cmd_valid_306), 
    .o_rdy(delay_stage_select[306] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_306), 
    .o_dat(tmp_icb_cmd_pack_306),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_307;
  wire     tmp_icb_cmd_valid_307;
  wire     tmp_icb_cmd_ready_307;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_307 (
    .i_vld(tmp_icb_cmd_valid_306), 
    .i_rdy(tmp_icb_cmd_ready_306), 
    .i_dat(tmp_icb_cmd_pack_306),
    .o_vld(tmp_icb_cmd_valid_307), 
    .o_rdy(delay_stage_select[307] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_307), 
    .o_dat(tmp_icb_cmd_pack_307),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_308;
  wire     tmp_icb_cmd_valid_308;
  wire     tmp_icb_cmd_ready_308;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_308 (
    .i_vld(tmp_icb_cmd_valid_307), 
    .i_rdy(tmp_icb_cmd_ready_307), 
    .i_dat(tmp_icb_cmd_pack_307),
    .o_vld(tmp_icb_cmd_valid_308), 
    .o_rdy(delay_stage_select[308] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_308), 
    .o_dat(tmp_icb_cmd_pack_308),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_309;
  wire     tmp_icb_cmd_valid_309;
  wire     tmp_icb_cmd_ready_309;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_309 (
    .i_vld(tmp_icb_cmd_valid_308), 
    .i_rdy(tmp_icb_cmd_ready_308), 
    .i_dat(tmp_icb_cmd_pack_308),
    .o_vld(tmp_icb_cmd_valid_309), 
    .o_rdy(delay_stage_select[309] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_309), 
    .o_dat(tmp_icb_cmd_pack_309),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_310;
  wire     tmp_icb_cmd_valid_310;
  wire     tmp_icb_cmd_ready_310;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_310 (
    .i_vld(tmp_icb_cmd_valid_309), 
    .i_rdy(tmp_icb_cmd_ready_309), 
    .i_dat(tmp_icb_cmd_pack_309),
    .o_vld(tmp_icb_cmd_valid_310), 
    .o_rdy(delay_stage_select[310] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_310), 
    .o_dat(tmp_icb_cmd_pack_310),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_311;
  wire     tmp_icb_cmd_valid_311;
  wire     tmp_icb_cmd_ready_311;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_311 (
    .i_vld(tmp_icb_cmd_valid_310), 
    .i_rdy(tmp_icb_cmd_ready_310), 
    .i_dat(tmp_icb_cmd_pack_310),
    .o_vld(tmp_icb_cmd_valid_311), 
    .o_rdy(delay_stage_select[311] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_311), 
    .o_dat(tmp_icb_cmd_pack_311),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_312;
  wire     tmp_icb_cmd_valid_312;
  wire     tmp_icb_cmd_ready_312;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_312 (
    .i_vld(tmp_icb_cmd_valid_311), 
    .i_rdy(tmp_icb_cmd_ready_311), 
    .i_dat(tmp_icb_cmd_pack_311),
    .o_vld(tmp_icb_cmd_valid_312), 
    .o_rdy(delay_stage_select[312] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_312), 
    .o_dat(tmp_icb_cmd_pack_312),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_313;
  wire     tmp_icb_cmd_valid_313;
  wire     tmp_icb_cmd_ready_313;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_313 (
    .i_vld(tmp_icb_cmd_valid_312), 
    .i_rdy(tmp_icb_cmd_ready_312), 
    .i_dat(tmp_icb_cmd_pack_312),
    .o_vld(tmp_icb_cmd_valid_313), 
    .o_rdy(delay_stage_select[313] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_313), 
    .o_dat(tmp_icb_cmd_pack_313),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_314;
  wire     tmp_icb_cmd_valid_314;
  wire     tmp_icb_cmd_ready_314;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_314 (
    .i_vld(tmp_icb_cmd_valid_313), 
    .i_rdy(tmp_icb_cmd_ready_313), 
    .i_dat(tmp_icb_cmd_pack_313),
    .o_vld(tmp_icb_cmd_valid_314), 
    .o_rdy(delay_stage_select[314] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_314), 
    .o_dat(tmp_icb_cmd_pack_314),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_315;
  wire     tmp_icb_cmd_valid_315;
  wire     tmp_icb_cmd_ready_315;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_315 (
    .i_vld(tmp_icb_cmd_valid_314), 
    .i_rdy(tmp_icb_cmd_ready_314), 
    .i_dat(tmp_icb_cmd_pack_314),
    .o_vld(tmp_icb_cmd_valid_315), 
    .o_rdy(delay_stage_select[315] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_315), 
    .o_dat(tmp_icb_cmd_pack_315),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_316;
  wire     tmp_icb_cmd_valid_316;
  wire     tmp_icb_cmd_ready_316;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_316 (
    .i_vld(tmp_icb_cmd_valid_315), 
    .i_rdy(tmp_icb_cmd_ready_315), 
    .i_dat(tmp_icb_cmd_pack_315),
    .o_vld(tmp_icb_cmd_valid_316), 
    .o_rdy(delay_stage_select[316] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_316), 
    .o_dat(tmp_icb_cmd_pack_316),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_317;
  wire     tmp_icb_cmd_valid_317;
  wire     tmp_icb_cmd_ready_317;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_317 (
    .i_vld(tmp_icb_cmd_valid_316), 
    .i_rdy(tmp_icb_cmd_ready_316), 
    .i_dat(tmp_icb_cmd_pack_316),
    .o_vld(tmp_icb_cmd_valid_317), 
    .o_rdy(delay_stage_select[317] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_317), 
    .o_dat(tmp_icb_cmd_pack_317),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_318;
  wire     tmp_icb_cmd_valid_318;
  wire     tmp_icb_cmd_ready_318;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_318 (
    .i_vld(tmp_icb_cmd_valid_317), 
    .i_rdy(tmp_icb_cmd_ready_317), 
    .i_dat(tmp_icb_cmd_pack_317),
    .o_vld(tmp_icb_cmd_valid_318), 
    .o_rdy(delay_stage_select[318] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_318), 
    .o_dat(tmp_icb_cmd_pack_318),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_319;
  wire     tmp_icb_cmd_valid_319;
  wire     tmp_icb_cmd_ready_319;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_319 (
    .i_vld(tmp_icb_cmd_valid_318), 
    .i_rdy(tmp_icb_cmd_ready_318), 
    .i_dat(tmp_icb_cmd_pack_318),
    .o_vld(tmp_icb_cmd_valid_319), 
    .o_rdy(delay_stage_select[319] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_319), 
    .o_dat(tmp_icb_cmd_pack_319),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_320;
  wire     tmp_icb_cmd_valid_320;
  wire     tmp_icb_cmd_ready_320;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_320 (
    .i_vld(tmp_icb_cmd_valid_319), 
    .i_rdy(tmp_icb_cmd_ready_319), 
    .i_dat(tmp_icb_cmd_pack_319),
    .o_vld(tmp_icb_cmd_valid_320), 
    .o_rdy(delay_stage_select[320] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_320), 
    .o_dat(tmp_icb_cmd_pack_320),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_321;
  wire     tmp_icb_cmd_valid_321;
  wire     tmp_icb_cmd_ready_321;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_321 (
    .i_vld(tmp_icb_cmd_valid_320), 
    .i_rdy(tmp_icb_cmd_ready_320), 
    .i_dat(tmp_icb_cmd_pack_320),
    .o_vld(tmp_icb_cmd_valid_321), 
    .o_rdy(delay_stage_select[321] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_321), 
    .o_dat(tmp_icb_cmd_pack_321),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_322;
  wire     tmp_icb_cmd_valid_322;
  wire     tmp_icb_cmd_ready_322;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_322 (
    .i_vld(tmp_icb_cmd_valid_321), 
    .i_rdy(tmp_icb_cmd_ready_321), 
    .i_dat(tmp_icb_cmd_pack_321),
    .o_vld(tmp_icb_cmd_valid_322), 
    .o_rdy(delay_stage_select[322] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_322), 
    .o_dat(tmp_icb_cmd_pack_322),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_323;
  wire     tmp_icb_cmd_valid_323;
  wire     tmp_icb_cmd_ready_323;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_323 (
    .i_vld(tmp_icb_cmd_valid_322), 
    .i_rdy(tmp_icb_cmd_ready_322), 
    .i_dat(tmp_icb_cmd_pack_322),
    .o_vld(tmp_icb_cmd_valid_323), 
    .o_rdy(delay_stage_select[323] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_323), 
    .o_dat(tmp_icb_cmd_pack_323),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_324;
  wire     tmp_icb_cmd_valid_324;
  wire     tmp_icb_cmd_ready_324;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_324 (
    .i_vld(tmp_icb_cmd_valid_323), 
    .i_rdy(tmp_icb_cmd_ready_323), 
    .i_dat(tmp_icb_cmd_pack_323),
    .o_vld(tmp_icb_cmd_valid_324), 
    .o_rdy(delay_stage_select[324] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_324), 
    .o_dat(tmp_icb_cmd_pack_324),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_325;
  wire     tmp_icb_cmd_valid_325;
  wire     tmp_icb_cmd_ready_325;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_325 (
    .i_vld(tmp_icb_cmd_valid_324), 
    .i_rdy(tmp_icb_cmd_ready_324), 
    .i_dat(tmp_icb_cmd_pack_324),
    .o_vld(tmp_icb_cmd_valid_325), 
    .o_rdy(delay_stage_select[325] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_325), 
    .o_dat(tmp_icb_cmd_pack_325),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_326;
  wire     tmp_icb_cmd_valid_326;
  wire     tmp_icb_cmd_ready_326;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_326 (
    .i_vld(tmp_icb_cmd_valid_325), 
    .i_rdy(tmp_icb_cmd_ready_325), 
    .i_dat(tmp_icb_cmd_pack_325),
    .o_vld(tmp_icb_cmd_valid_326), 
    .o_rdy(delay_stage_select[326] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_326), 
    .o_dat(tmp_icb_cmd_pack_326),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_327;
  wire     tmp_icb_cmd_valid_327;
  wire     tmp_icb_cmd_ready_327;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_327 (
    .i_vld(tmp_icb_cmd_valid_326), 
    .i_rdy(tmp_icb_cmd_ready_326), 
    .i_dat(tmp_icb_cmd_pack_326),
    .o_vld(tmp_icb_cmd_valid_327), 
    .o_rdy(delay_stage_select[327] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_327), 
    .o_dat(tmp_icb_cmd_pack_327),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_328;
  wire     tmp_icb_cmd_valid_328;
  wire     tmp_icb_cmd_ready_328;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_328 (
    .i_vld(tmp_icb_cmd_valid_327), 
    .i_rdy(tmp_icb_cmd_ready_327), 
    .i_dat(tmp_icb_cmd_pack_327),
    .o_vld(tmp_icb_cmd_valid_328), 
    .o_rdy(delay_stage_select[328] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_328), 
    .o_dat(tmp_icb_cmd_pack_328),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_329;
  wire     tmp_icb_cmd_valid_329;
  wire     tmp_icb_cmd_ready_329;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_329 (
    .i_vld(tmp_icb_cmd_valid_328), 
    .i_rdy(tmp_icb_cmd_ready_328), 
    .i_dat(tmp_icb_cmd_pack_328),
    .o_vld(tmp_icb_cmd_valid_329), 
    .o_rdy(delay_stage_select[329] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_329), 
    .o_dat(tmp_icb_cmd_pack_329),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_330;
  wire     tmp_icb_cmd_valid_330;
  wire     tmp_icb_cmd_ready_330;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_330 (
    .i_vld(tmp_icb_cmd_valid_329), 
    .i_rdy(tmp_icb_cmd_ready_329), 
    .i_dat(tmp_icb_cmd_pack_329),
    .o_vld(tmp_icb_cmd_valid_330), 
    .o_rdy(delay_stage_select[330] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_330), 
    .o_dat(tmp_icb_cmd_pack_330),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_331;
  wire     tmp_icb_cmd_valid_331;
  wire     tmp_icb_cmd_ready_331;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_331 (
    .i_vld(tmp_icb_cmd_valid_330), 
    .i_rdy(tmp_icb_cmd_ready_330), 
    .i_dat(tmp_icb_cmd_pack_330),
    .o_vld(tmp_icb_cmd_valid_331), 
    .o_rdy(delay_stage_select[331] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_331), 
    .o_dat(tmp_icb_cmd_pack_331),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_332;
  wire     tmp_icb_cmd_valid_332;
  wire     tmp_icb_cmd_ready_332;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_332 (
    .i_vld(tmp_icb_cmd_valid_331), 
    .i_rdy(tmp_icb_cmd_ready_331), 
    .i_dat(tmp_icb_cmd_pack_331),
    .o_vld(tmp_icb_cmd_valid_332), 
    .o_rdy(delay_stage_select[332] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_332), 
    .o_dat(tmp_icb_cmd_pack_332),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_333;
  wire     tmp_icb_cmd_valid_333;
  wire     tmp_icb_cmd_ready_333;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_333 (
    .i_vld(tmp_icb_cmd_valid_332), 
    .i_rdy(tmp_icb_cmd_ready_332), 
    .i_dat(tmp_icb_cmd_pack_332),
    .o_vld(tmp_icb_cmd_valid_333), 
    .o_rdy(delay_stage_select[333] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_333), 
    .o_dat(tmp_icb_cmd_pack_333),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_334;
  wire     tmp_icb_cmd_valid_334;
  wire     tmp_icb_cmd_ready_334;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_334 (
    .i_vld(tmp_icb_cmd_valid_333), 
    .i_rdy(tmp_icb_cmd_ready_333), 
    .i_dat(tmp_icb_cmd_pack_333),
    .o_vld(tmp_icb_cmd_valid_334), 
    .o_rdy(delay_stage_select[334] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_334), 
    .o_dat(tmp_icb_cmd_pack_334),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_335;
  wire     tmp_icb_cmd_valid_335;
  wire     tmp_icb_cmd_ready_335;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_335 (
    .i_vld(tmp_icb_cmd_valid_334), 
    .i_rdy(tmp_icb_cmd_ready_334), 
    .i_dat(tmp_icb_cmd_pack_334),
    .o_vld(tmp_icb_cmd_valid_335), 
    .o_rdy(delay_stage_select[335] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_335), 
    .o_dat(tmp_icb_cmd_pack_335),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_336;
  wire     tmp_icb_cmd_valid_336;
  wire     tmp_icb_cmd_ready_336;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_336 (
    .i_vld(tmp_icb_cmd_valid_335), 
    .i_rdy(tmp_icb_cmd_ready_335), 
    .i_dat(tmp_icb_cmd_pack_335),
    .o_vld(tmp_icb_cmd_valid_336), 
    .o_rdy(delay_stage_select[336] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_336), 
    .o_dat(tmp_icb_cmd_pack_336),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_337;
  wire     tmp_icb_cmd_valid_337;
  wire     tmp_icb_cmd_ready_337;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_337 (
    .i_vld(tmp_icb_cmd_valid_336), 
    .i_rdy(tmp_icb_cmd_ready_336), 
    .i_dat(tmp_icb_cmd_pack_336),
    .o_vld(tmp_icb_cmd_valid_337), 
    .o_rdy(delay_stage_select[337] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_337), 
    .o_dat(tmp_icb_cmd_pack_337),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_338;
  wire     tmp_icb_cmd_valid_338;
  wire     tmp_icb_cmd_ready_338;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_338 (
    .i_vld(tmp_icb_cmd_valid_337), 
    .i_rdy(tmp_icb_cmd_ready_337), 
    .i_dat(tmp_icb_cmd_pack_337),
    .o_vld(tmp_icb_cmd_valid_338), 
    .o_rdy(delay_stage_select[338] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_338), 
    .o_dat(tmp_icb_cmd_pack_338),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_339;
  wire     tmp_icb_cmd_valid_339;
  wire     tmp_icb_cmd_ready_339;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_339 (
    .i_vld(tmp_icb_cmd_valid_338), 
    .i_rdy(tmp_icb_cmd_ready_338), 
    .i_dat(tmp_icb_cmd_pack_338),
    .o_vld(tmp_icb_cmd_valid_339), 
    .o_rdy(delay_stage_select[339] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_339), 
    .o_dat(tmp_icb_cmd_pack_339),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_340;
  wire     tmp_icb_cmd_valid_340;
  wire     tmp_icb_cmd_ready_340;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_340 (
    .i_vld(tmp_icb_cmd_valid_339), 
    .i_rdy(tmp_icb_cmd_ready_339), 
    .i_dat(tmp_icb_cmd_pack_339),
    .o_vld(tmp_icb_cmd_valid_340), 
    .o_rdy(delay_stage_select[340] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_340), 
    .o_dat(tmp_icb_cmd_pack_340),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_341;
  wire     tmp_icb_cmd_valid_341;
  wire     tmp_icb_cmd_ready_341;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_341 (
    .i_vld(tmp_icb_cmd_valid_340), 
    .i_rdy(tmp_icb_cmd_ready_340), 
    .i_dat(tmp_icb_cmd_pack_340),
    .o_vld(tmp_icb_cmd_valid_341), 
    .o_rdy(delay_stage_select[341] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_341), 
    .o_dat(tmp_icb_cmd_pack_341),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_342;
  wire     tmp_icb_cmd_valid_342;
  wire     tmp_icb_cmd_ready_342;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_342 (
    .i_vld(tmp_icb_cmd_valid_341), 
    .i_rdy(tmp_icb_cmd_ready_341), 
    .i_dat(tmp_icb_cmd_pack_341),
    .o_vld(tmp_icb_cmd_valid_342), 
    .o_rdy(delay_stage_select[342] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_342), 
    .o_dat(tmp_icb_cmd_pack_342),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_343;
  wire     tmp_icb_cmd_valid_343;
  wire     tmp_icb_cmd_ready_343;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_343 (
    .i_vld(tmp_icb_cmd_valid_342), 
    .i_rdy(tmp_icb_cmd_ready_342), 
    .i_dat(tmp_icb_cmd_pack_342),
    .o_vld(tmp_icb_cmd_valid_343), 
    .o_rdy(delay_stage_select[343] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_343), 
    .o_dat(tmp_icb_cmd_pack_343),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_344;
  wire     tmp_icb_cmd_valid_344;
  wire     tmp_icb_cmd_ready_344;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_344 (
    .i_vld(tmp_icb_cmd_valid_343), 
    .i_rdy(tmp_icb_cmd_ready_343), 
    .i_dat(tmp_icb_cmd_pack_343),
    .o_vld(tmp_icb_cmd_valid_344), 
    .o_rdy(delay_stage_select[344] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_344), 
    .o_dat(tmp_icb_cmd_pack_344),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_345;
  wire     tmp_icb_cmd_valid_345;
  wire     tmp_icb_cmd_ready_345;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_345 (
    .i_vld(tmp_icb_cmd_valid_344), 
    .i_rdy(tmp_icb_cmd_ready_344), 
    .i_dat(tmp_icb_cmd_pack_344),
    .o_vld(tmp_icb_cmd_valid_345), 
    .o_rdy(delay_stage_select[345] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_345), 
    .o_dat(tmp_icb_cmd_pack_345),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_346;
  wire     tmp_icb_cmd_valid_346;
  wire     tmp_icb_cmd_ready_346;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_346 (
    .i_vld(tmp_icb_cmd_valid_345), 
    .i_rdy(tmp_icb_cmd_ready_345), 
    .i_dat(tmp_icb_cmd_pack_345),
    .o_vld(tmp_icb_cmd_valid_346), 
    .o_rdy(delay_stage_select[346] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_346), 
    .o_dat(tmp_icb_cmd_pack_346),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_347;
  wire     tmp_icb_cmd_valid_347;
  wire     tmp_icb_cmd_ready_347;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_347 (
    .i_vld(tmp_icb_cmd_valid_346), 
    .i_rdy(tmp_icb_cmd_ready_346), 
    .i_dat(tmp_icb_cmd_pack_346),
    .o_vld(tmp_icb_cmd_valid_347), 
    .o_rdy(delay_stage_select[347] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_347), 
    .o_dat(tmp_icb_cmd_pack_347),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_348;
  wire     tmp_icb_cmd_valid_348;
  wire     tmp_icb_cmd_ready_348;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_348 (
    .i_vld(tmp_icb_cmd_valid_347), 
    .i_rdy(tmp_icb_cmd_ready_347), 
    .i_dat(tmp_icb_cmd_pack_347),
    .o_vld(tmp_icb_cmd_valid_348), 
    .o_rdy(delay_stage_select[348] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_348), 
    .o_dat(tmp_icb_cmd_pack_348),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_349;
  wire     tmp_icb_cmd_valid_349;
  wire     tmp_icb_cmd_ready_349;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_349 (
    .i_vld(tmp_icb_cmd_valid_348), 
    .i_rdy(tmp_icb_cmd_ready_348), 
    .i_dat(tmp_icb_cmd_pack_348),
    .o_vld(tmp_icb_cmd_valid_349), 
    .o_rdy(delay_stage_select[349] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_349), 
    .o_dat(tmp_icb_cmd_pack_349),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_350;
  wire     tmp_icb_cmd_valid_350;
  wire     tmp_icb_cmd_ready_350;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_350 (
    .i_vld(tmp_icb_cmd_valid_349), 
    .i_rdy(tmp_icb_cmd_ready_349), 
    .i_dat(tmp_icb_cmd_pack_349),
    .o_vld(tmp_icb_cmd_valid_350), 
    .o_rdy(delay_stage_select[350] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_350), 
    .o_dat(tmp_icb_cmd_pack_350),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_351;
  wire     tmp_icb_cmd_valid_351;
  wire     tmp_icb_cmd_ready_351;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_351 (
    .i_vld(tmp_icb_cmd_valid_350), 
    .i_rdy(tmp_icb_cmd_ready_350), 
    .i_dat(tmp_icb_cmd_pack_350),
    .o_vld(tmp_icb_cmd_valid_351), 
    .o_rdy(delay_stage_select[351] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_351), 
    .o_dat(tmp_icb_cmd_pack_351),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_352;
  wire     tmp_icb_cmd_valid_352;
  wire     tmp_icb_cmd_ready_352;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_352 (
    .i_vld(tmp_icb_cmd_valid_351), 
    .i_rdy(tmp_icb_cmd_ready_351), 
    .i_dat(tmp_icb_cmd_pack_351),
    .o_vld(tmp_icb_cmd_valid_352), 
    .o_rdy(delay_stage_select[352] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_352), 
    .o_dat(tmp_icb_cmd_pack_352),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_353;
  wire     tmp_icb_cmd_valid_353;
  wire     tmp_icb_cmd_ready_353;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_353 (
    .i_vld(tmp_icb_cmd_valid_352), 
    .i_rdy(tmp_icb_cmd_ready_352), 
    .i_dat(tmp_icb_cmd_pack_352),
    .o_vld(tmp_icb_cmd_valid_353), 
    .o_rdy(delay_stage_select[353] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_353), 
    .o_dat(tmp_icb_cmd_pack_353),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_354;
  wire     tmp_icb_cmd_valid_354;
  wire     tmp_icb_cmd_ready_354;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_354 (
    .i_vld(tmp_icb_cmd_valid_353), 
    .i_rdy(tmp_icb_cmd_ready_353), 
    .i_dat(tmp_icb_cmd_pack_353),
    .o_vld(tmp_icb_cmd_valid_354), 
    .o_rdy(delay_stage_select[354] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_354), 
    .o_dat(tmp_icb_cmd_pack_354),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_355;
  wire     tmp_icb_cmd_valid_355;
  wire     tmp_icb_cmd_ready_355;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_355 (
    .i_vld(tmp_icb_cmd_valid_354), 
    .i_rdy(tmp_icb_cmd_ready_354), 
    .i_dat(tmp_icb_cmd_pack_354),
    .o_vld(tmp_icb_cmd_valid_355), 
    .o_rdy(delay_stage_select[355] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_355), 
    .o_dat(tmp_icb_cmd_pack_355),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_356;
  wire     tmp_icb_cmd_valid_356;
  wire     tmp_icb_cmd_ready_356;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_356 (
    .i_vld(tmp_icb_cmd_valid_355), 
    .i_rdy(tmp_icb_cmd_ready_355), 
    .i_dat(tmp_icb_cmd_pack_355),
    .o_vld(tmp_icb_cmd_valid_356), 
    .o_rdy(delay_stage_select[356] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_356), 
    .o_dat(tmp_icb_cmd_pack_356),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_357;
  wire     tmp_icb_cmd_valid_357;
  wire     tmp_icb_cmd_ready_357;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_357 (
    .i_vld(tmp_icb_cmd_valid_356), 
    .i_rdy(tmp_icb_cmd_ready_356), 
    .i_dat(tmp_icb_cmd_pack_356),
    .o_vld(tmp_icb_cmd_valid_357), 
    .o_rdy(delay_stage_select[357] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_357), 
    .o_dat(tmp_icb_cmd_pack_357),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_358;
  wire     tmp_icb_cmd_valid_358;
  wire     tmp_icb_cmd_ready_358;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_358 (
    .i_vld(tmp_icb_cmd_valid_357), 
    .i_rdy(tmp_icb_cmd_ready_357), 
    .i_dat(tmp_icb_cmd_pack_357),
    .o_vld(tmp_icb_cmd_valid_358), 
    .o_rdy(delay_stage_select[358] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_358), 
    .o_dat(tmp_icb_cmd_pack_358),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_359;
  wire     tmp_icb_cmd_valid_359;
  wire     tmp_icb_cmd_ready_359;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_359 (
    .i_vld(tmp_icb_cmd_valid_358), 
    .i_rdy(tmp_icb_cmd_ready_358), 
    .i_dat(tmp_icb_cmd_pack_358),
    .o_vld(tmp_icb_cmd_valid_359), 
    .o_rdy(delay_stage_select[359] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_359), 
    .o_dat(tmp_icb_cmd_pack_359),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_360;
  wire     tmp_icb_cmd_valid_360;
  wire     tmp_icb_cmd_ready_360;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_360 (
    .i_vld(tmp_icb_cmd_valid_359), 
    .i_rdy(tmp_icb_cmd_ready_359), 
    .i_dat(tmp_icb_cmd_pack_359),
    .o_vld(tmp_icb_cmd_valid_360), 
    .o_rdy(delay_stage_select[360] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_360), 
    .o_dat(tmp_icb_cmd_pack_360),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_361;
  wire     tmp_icb_cmd_valid_361;
  wire     tmp_icb_cmd_ready_361;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_361 (
    .i_vld(tmp_icb_cmd_valid_360), 
    .i_rdy(tmp_icb_cmd_ready_360), 
    .i_dat(tmp_icb_cmd_pack_360),
    .o_vld(tmp_icb_cmd_valid_361), 
    .o_rdy(delay_stage_select[361] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_361), 
    .o_dat(tmp_icb_cmd_pack_361),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_362;
  wire     tmp_icb_cmd_valid_362;
  wire     tmp_icb_cmd_ready_362;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_362 (
    .i_vld(tmp_icb_cmd_valid_361), 
    .i_rdy(tmp_icb_cmd_ready_361), 
    .i_dat(tmp_icb_cmd_pack_361),
    .o_vld(tmp_icb_cmd_valid_362), 
    .o_rdy(delay_stage_select[362] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_362), 
    .o_dat(tmp_icb_cmd_pack_362),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_363;
  wire     tmp_icb_cmd_valid_363;
  wire     tmp_icb_cmd_ready_363;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_363 (
    .i_vld(tmp_icb_cmd_valid_362), 
    .i_rdy(tmp_icb_cmd_ready_362), 
    .i_dat(tmp_icb_cmd_pack_362),
    .o_vld(tmp_icb_cmd_valid_363), 
    .o_rdy(delay_stage_select[363] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_363), 
    .o_dat(tmp_icb_cmd_pack_363),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_364;
  wire     tmp_icb_cmd_valid_364;
  wire     tmp_icb_cmd_ready_364;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_364 (
    .i_vld(tmp_icb_cmd_valid_363), 
    .i_rdy(tmp_icb_cmd_ready_363), 
    .i_dat(tmp_icb_cmd_pack_363),
    .o_vld(tmp_icb_cmd_valid_364), 
    .o_rdy(delay_stage_select[364] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_364), 
    .o_dat(tmp_icb_cmd_pack_364),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_365;
  wire     tmp_icb_cmd_valid_365;
  wire     tmp_icb_cmd_ready_365;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_365 (
    .i_vld(tmp_icb_cmd_valid_364), 
    .i_rdy(tmp_icb_cmd_ready_364), 
    .i_dat(tmp_icb_cmd_pack_364),
    .o_vld(tmp_icb_cmd_valid_365), 
    .o_rdy(delay_stage_select[365] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_365), 
    .o_dat(tmp_icb_cmd_pack_365),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_366;
  wire     tmp_icb_cmd_valid_366;
  wire     tmp_icb_cmd_ready_366;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_366 (
    .i_vld(tmp_icb_cmd_valid_365), 
    .i_rdy(tmp_icb_cmd_ready_365), 
    .i_dat(tmp_icb_cmd_pack_365),
    .o_vld(tmp_icb_cmd_valid_366), 
    .o_rdy(delay_stage_select[366] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_366), 
    .o_dat(tmp_icb_cmd_pack_366),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_367;
  wire     tmp_icb_cmd_valid_367;
  wire     tmp_icb_cmd_ready_367;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_367 (
    .i_vld(tmp_icb_cmd_valid_366), 
    .i_rdy(tmp_icb_cmd_ready_366), 
    .i_dat(tmp_icb_cmd_pack_366),
    .o_vld(tmp_icb_cmd_valid_367), 
    .o_rdy(delay_stage_select[367] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_367), 
    .o_dat(tmp_icb_cmd_pack_367),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_368;
  wire     tmp_icb_cmd_valid_368;
  wire     tmp_icb_cmd_ready_368;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_368 (
    .i_vld(tmp_icb_cmd_valid_367), 
    .i_rdy(tmp_icb_cmd_ready_367), 
    .i_dat(tmp_icb_cmd_pack_367),
    .o_vld(tmp_icb_cmd_valid_368), 
    .o_rdy(delay_stage_select[368] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_368), 
    .o_dat(tmp_icb_cmd_pack_368),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_369;
  wire     tmp_icb_cmd_valid_369;
  wire     tmp_icb_cmd_ready_369;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_369 (
    .i_vld(tmp_icb_cmd_valid_368), 
    .i_rdy(tmp_icb_cmd_ready_368), 
    .i_dat(tmp_icb_cmd_pack_368),
    .o_vld(tmp_icb_cmd_valid_369), 
    .o_rdy(delay_stage_select[369] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_369), 
    .o_dat(tmp_icb_cmd_pack_369),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_370;
  wire     tmp_icb_cmd_valid_370;
  wire     tmp_icb_cmd_ready_370;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_370 (
    .i_vld(tmp_icb_cmd_valid_369), 
    .i_rdy(tmp_icb_cmd_ready_369), 
    .i_dat(tmp_icb_cmd_pack_369),
    .o_vld(tmp_icb_cmd_valid_370), 
    .o_rdy(delay_stage_select[370] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_370), 
    .o_dat(tmp_icb_cmd_pack_370),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_371;
  wire     tmp_icb_cmd_valid_371;
  wire     tmp_icb_cmd_ready_371;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_371 (
    .i_vld(tmp_icb_cmd_valid_370), 
    .i_rdy(tmp_icb_cmd_ready_370), 
    .i_dat(tmp_icb_cmd_pack_370),
    .o_vld(tmp_icb_cmd_valid_371), 
    .o_rdy(delay_stage_select[371] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_371), 
    .o_dat(tmp_icb_cmd_pack_371),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_372;
  wire     tmp_icb_cmd_valid_372;
  wire     tmp_icb_cmd_ready_372;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_372 (
    .i_vld(tmp_icb_cmd_valid_371), 
    .i_rdy(tmp_icb_cmd_ready_371), 
    .i_dat(tmp_icb_cmd_pack_371),
    .o_vld(tmp_icb_cmd_valid_372), 
    .o_rdy(delay_stage_select[372] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_372), 
    .o_dat(tmp_icb_cmd_pack_372),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_373;
  wire     tmp_icb_cmd_valid_373;
  wire     tmp_icb_cmd_ready_373;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_373 (
    .i_vld(tmp_icb_cmd_valid_372), 
    .i_rdy(tmp_icb_cmd_ready_372), 
    .i_dat(tmp_icb_cmd_pack_372),
    .o_vld(tmp_icb_cmd_valid_373), 
    .o_rdy(delay_stage_select[373] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_373), 
    .o_dat(tmp_icb_cmd_pack_373),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_374;
  wire     tmp_icb_cmd_valid_374;
  wire     tmp_icb_cmd_ready_374;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_374 (
    .i_vld(tmp_icb_cmd_valid_373), 
    .i_rdy(tmp_icb_cmd_ready_373), 
    .i_dat(tmp_icb_cmd_pack_373),
    .o_vld(tmp_icb_cmd_valid_374), 
    .o_rdy(delay_stage_select[374] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_374), 
    .o_dat(tmp_icb_cmd_pack_374),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_375;
  wire     tmp_icb_cmd_valid_375;
  wire     tmp_icb_cmd_ready_375;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_375 (
    .i_vld(tmp_icb_cmd_valid_374), 
    .i_rdy(tmp_icb_cmd_ready_374), 
    .i_dat(tmp_icb_cmd_pack_374),
    .o_vld(tmp_icb_cmd_valid_375), 
    .o_rdy(delay_stage_select[375] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_375), 
    .o_dat(tmp_icb_cmd_pack_375),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_376;
  wire     tmp_icb_cmd_valid_376;
  wire     tmp_icb_cmd_ready_376;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_376 (
    .i_vld(tmp_icb_cmd_valid_375), 
    .i_rdy(tmp_icb_cmd_ready_375), 
    .i_dat(tmp_icb_cmd_pack_375),
    .o_vld(tmp_icb_cmd_valid_376), 
    .o_rdy(delay_stage_select[376] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_376), 
    .o_dat(tmp_icb_cmd_pack_376),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_377;
  wire     tmp_icb_cmd_valid_377;
  wire     tmp_icb_cmd_ready_377;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_377 (
    .i_vld(tmp_icb_cmd_valid_376), 
    .i_rdy(tmp_icb_cmd_ready_376), 
    .i_dat(tmp_icb_cmd_pack_376),
    .o_vld(tmp_icb_cmd_valid_377), 
    .o_rdy(delay_stage_select[377] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_377), 
    .o_dat(tmp_icb_cmd_pack_377),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_378;
  wire     tmp_icb_cmd_valid_378;
  wire     tmp_icb_cmd_ready_378;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_378 (
    .i_vld(tmp_icb_cmd_valid_377), 
    .i_rdy(tmp_icb_cmd_ready_377), 
    .i_dat(tmp_icb_cmd_pack_377),
    .o_vld(tmp_icb_cmd_valid_378), 
    .o_rdy(delay_stage_select[378] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_378), 
    .o_dat(tmp_icb_cmd_pack_378),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_379;
  wire     tmp_icb_cmd_valid_379;
  wire     tmp_icb_cmd_ready_379;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_379 (
    .i_vld(tmp_icb_cmd_valid_378), 
    .i_rdy(tmp_icb_cmd_ready_378), 
    .i_dat(tmp_icb_cmd_pack_378),
    .o_vld(tmp_icb_cmd_valid_379), 
    .o_rdy(delay_stage_select[379] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_379), 
    .o_dat(tmp_icb_cmd_pack_379),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_380;
  wire     tmp_icb_cmd_valid_380;
  wire     tmp_icb_cmd_ready_380;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_380 (
    .i_vld(tmp_icb_cmd_valid_379), 
    .i_rdy(tmp_icb_cmd_ready_379), 
    .i_dat(tmp_icb_cmd_pack_379),
    .o_vld(tmp_icb_cmd_valid_380), 
    .o_rdy(delay_stage_select[380] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_380), 
    .o_dat(tmp_icb_cmd_pack_380),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_381;
  wire     tmp_icb_cmd_valid_381;
  wire     tmp_icb_cmd_ready_381;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_381 (
    .i_vld(tmp_icb_cmd_valid_380), 
    .i_rdy(tmp_icb_cmd_ready_380), 
    .i_dat(tmp_icb_cmd_pack_380),
    .o_vld(tmp_icb_cmd_valid_381), 
    .o_rdy(delay_stage_select[381] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_381), 
    .o_dat(tmp_icb_cmd_pack_381),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_382;
  wire     tmp_icb_cmd_valid_382;
  wire     tmp_icb_cmd_ready_382;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_382 (
    .i_vld(tmp_icb_cmd_valid_381), 
    .i_rdy(tmp_icb_cmd_ready_381), 
    .i_dat(tmp_icb_cmd_pack_381),
    .o_vld(tmp_icb_cmd_valid_382), 
    .o_rdy(delay_stage_select[382] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_382), 
    .o_dat(tmp_icb_cmd_pack_382),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_383;
  wire     tmp_icb_cmd_valid_383;
  wire     tmp_icb_cmd_ready_383;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_383 (
    .i_vld(tmp_icb_cmd_valid_382), 
    .i_rdy(tmp_icb_cmd_ready_382), 
    .i_dat(tmp_icb_cmd_pack_382),
    .o_vld(tmp_icb_cmd_valid_383), 
    .o_rdy(delay_stage_select[383] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_383), 
    .o_dat(tmp_icb_cmd_pack_383),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_384;
  wire     tmp_icb_cmd_valid_384;
  wire     tmp_icb_cmd_ready_384;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_384 (
    .i_vld(tmp_icb_cmd_valid_383), 
    .i_rdy(tmp_icb_cmd_ready_383), 
    .i_dat(tmp_icb_cmd_pack_383),
    .o_vld(tmp_icb_cmd_valid_384), 
    .o_rdy(delay_stage_select[384] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_384), 
    .o_dat(tmp_icb_cmd_pack_384),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_385;
  wire     tmp_icb_cmd_valid_385;
  wire     tmp_icb_cmd_ready_385;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_385 (
    .i_vld(tmp_icb_cmd_valid_384), 
    .i_rdy(tmp_icb_cmd_ready_384), 
    .i_dat(tmp_icb_cmd_pack_384),
    .o_vld(tmp_icb_cmd_valid_385), 
    .o_rdy(delay_stage_select[385] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_385), 
    .o_dat(tmp_icb_cmd_pack_385),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_386;
  wire     tmp_icb_cmd_valid_386;
  wire     tmp_icb_cmd_ready_386;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_386 (
    .i_vld(tmp_icb_cmd_valid_385), 
    .i_rdy(tmp_icb_cmd_ready_385), 
    .i_dat(tmp_icb_cmd_pack_385),
    .o_vld(tmp_icb_cmd_valid_386), 
    .o_rdy(delay_stage_select[386] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_386), 
    .o_dat(tmp_icb_cmd_pack_386),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_387;
  wire     tmp_icb_cmd_valid_387;
  wire     tmp_icb_cmd_ready_387;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_387 (
    .i_vld(tmp_icb_cmd_valid_386), 
    .i_rdy(tmp_icb_cmd_ready_386), 
    .i_dat(tmp_icb_cmd_pack_386),
    .o_vld(tmp_icb_cmd_valid_387), 
    .o_rdy(delay_stage_select[387] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_387), 
    .o_dat(tmp_icb_cmd_pack_387),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_388;
  wire     tmp_icb_cmd_valid_388;
  wire     tmp_icb_cmd_ready_388;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_388 (
    .i_vld(tmp_icb_cmd_valid_387), 
    .i_rdy(tmp_icb_cmd_ready_387), 
    .i_dat(tmp_icb_cmd_pack_387),
    .o_vld(tmp_icb_cmd_valid_388), 
    .o_rdy(delay_stage_select[388] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_388), 
    .o_dat(tmp_icb_cmd_pack_388),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_389;
  wire     tmp_icb_cmd_valid_389;
  wire     tmp_icb_cmd_ready_389;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_389 (
    .i_vld(tmp_icb_cmd_valid_388), 
    .i_rdy(tmp_icb_cmd_ready_388), 
    .i_dat(tmp_icb_cmd_pack_388),
    .o_vld(tmp_icb_cmd_valid_389), 
    .o_rdy(delay_stage_select[389] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_389), 
    .o_dat(tmp_icb_cmd_pack_389),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_390;
  wire     tmp_icb_cmd_valid_390;
  wire     tmp_icb_cmd_ready_390;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_390 (
    .i_vld(tmp_icb_cmd_valid_389), 
    .i_rdy(tmp_icb_cmd_ready_389), 
    .i_dat(tmp_icb_cmd_pack_389),
    .o_vld(tmp_icb_cmd_valid_390), 
    .o_rdy(delay_stage_select[390] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_390), 
    .o_dat(tmp_icb_cmd_pack_390),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_391;
  wire     tmp_icb_cmd_valid_391;
  wire     tmp_icb_cmd_ready_391;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_391 (
    .i_vld(tmp_icb_cmd_valid_390), 
    .i_rdy(tmp_icb_cmd_ready_390), 
    .i_dat(tmp_icb_cmd_pack_390),
    .o_vld(tmp_icb_cmd_valid_391), 
    .o_rdy(delay_stage_select[391] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_391), 
    .o_dat(tmp_icb_cmd_pack_391),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_392;
  wire     tmp_icb_cmd_valid_392;
  wire     tmp_icb_cmd_ready_392;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_392 (
    .i_vld(tmp_icb_cmd_valid_391), 
    .i_rdy(tmp_icb_cmd_ready_391), 
    .i_dat(tmp_icb_cmd_pack_391),
    .o_vld(tmp_icb_cmd_valid_392), 
    .o_rdy(delay_stage_select[392] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_392), 
    .o_dat(tmp_icb_cmd_pack_392),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_393;
  wire     tmp_icb_cmd_valid_393;
  wire     tmp_icb_cmd_ready_393;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_393 (
    .i_vld(tmp_icb_cmd_valid_392), 
    .i_rdy(tmp_icb_cmd_ready_392), 
    .i_dat(tmp_icb_cmd_pack_392),
    .o_vld(tmp_icb_cmd_valid_393), 
    .o_rdy(delay_stage_select[393] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_393), 
    .o_dat(tmp_icb_cmd_pack_393),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_394;
  wire     tmp_icb_cmd_valid_394;
  wire     tmp_icb_cmd_ready_394;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_394 (
    .i_vld(tmp_icb_cmd_valid_393), 
    .i_rdy(tmp_icb_cmd_ready_393), 
    .i_dat(tmp_icb_cmd_pack_393),
    .o_vld(tmp_icb_cmd_valid_394), 
    .o_rdy(delay_stage_select[394] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_394), 
    .o_dat(tmp_icb_cmd_pack_394),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_395;
  wire     tmp_icb_cmd_valid_395;
  wire     tmp_icb_cmd_ready_395;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_395 (
    .i_vld(tmp_icb_cmd_valid_394), 
    .i_rdy(tmp_icb_cmd_ready_394), 
    .i_dat(tmp_icb_cmd_pack_394),
    .o_vld(tmp_icb_cmd_valid_395), 
    .o_rdy(delay_stage_select[395] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_395), 
    .o_dat(tmp_icb_cmd_pack_395),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_396;
  wire     tmp_icb_cmd_valid_396;
  wire     tmp_icb_cmd_ready_396;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_396 (
    .i_vld(tmp_icb_cmd_valid_395), 
    .i_rdy(tmp_icb_cmd_ready_395), 
    .i_dat(tmp_icb_cmd_pack_395),
    .o_vld(tmp_icb_cmd_valid_396), 
    .o_rdy(delay_stage_select[396] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_396), 
    .o_dat(tmp_icb_cmd_pack_396),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_397;
  wire     tmp_icb_cmd_valid_397;
  wire     tmp_icb_cmd_ready_397;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_397 (
    .i_vld(tmp_icb_cmd_valid_396), 
    .i_rdy(tmp_icb_cmd_ready_396), 
    .i_dat(tmp_icb_cmd_pack_396),
    .o_vld(tmp_icb_cmd_valid_397), 
    .o_rdy(delay_stage_select[397] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_397), 
    .o_dat(tmp_icb_cmd_pack_397),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_398;
  wire     tmp_icb_cmd_valid_398;
  wire     tmp_icb_cmd_ready_398;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_398 (
    .i_vld(tmp_icb_cmd_valid_397), 
    .i_rdy(tmp_icb_cmd_ready_397), 
    .i_dat(tmp_icb_cmd_pack_397),
    .o_vld(tmp_icb_cmd_valid_398), 
    .o_rdy(delay_stage_select[398] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_398), 
    .o_dat(tmp_icb_cmd_pack_398),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_399;
  wire     tmp_icb_cmd_valid_399;
  wire     tmp_icb_cmd_ready_399;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_399 (
    .i_vld(tmp_icb_cmd_valid_398), 
    .i_rdy(tmp_icb_cmd_ready_398), 
    .i_dat(tmp_icb_cmd_pack_398),
    .o_vld(tmp_icb_cmd_valid_399), 
    .o_rdy(delay_stage_select[399] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_399), 
    .o_dat(tmp_icb_cmd_pack_399),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_400;
  wire     tmp_icb_cmd_valid_400;
  wire     tmp_icb_cmd_ready_400;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_400 (
    .i_vld(tmp_icb_cmd_valid_399), 
    .i_rdy(tmp_icb_cmd_ready_399), 
    .i_dat(tmp_icb_cmd_pack_399),
    .o_vld(tmp_icb_cmd_valid_400), 
    .o_rdy(delay_stage_select[400] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_400), 
    .o_dat(tmp_icb_cmd_pack_400),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_401;
  wire     tmp_icb_cmd_valid_401;
  wire     tmp_icb_cmd_ready_401;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_401 (
    .i_vld(tmp_icb_cmd_valid_400), 
    .i_rdy(tmp_icb_cmd_ready_400), 
    .i_dat(tmp_icb_cmd_pack_400),
    .o_vld(tmp_icb_cmd_valid_401), 
    .o_rdy(delay_stage_select[401] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_401), 
    .o_dat(tmp_icb_cmd_pack_401),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_402;
  wire     tmp_icb_cmd_valid_402;
  wire     tmp_icb_cmd_ready_402;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_402 (
    .i_vld(tmp_icb_cmd_valid_401), 
    .i_rdy(tmp_icb_cmd_ready_401), 
    .i_dat(tmp_icb_cmd_pack_401),
    .o_vld(tmp_icb_cmd_valid_402), 
    .o_rdy(delay_stage_select[402] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_402), 
    .o_dat(tmp_icb_cmd_pack_402),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_403;
  wire     tmp_icb_cmd_valid_403;
  wire     tmp_icb_cmd_ready_403;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_403 (
    .i_vld(tmp_icb_cmd_valid_402), 
    .i_rdy(tmp_icb_cmd_ready_402), 
    .i_dat(tmp_icb_cmd_pack_402),
    .o_vld(tmp_icb_cmd_valid_403), 
    .o_rdy(delay_stage_select[403] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_403), 
    .o_dat(tmp_icb_cmd_pack_403),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_404;
  wire     tmp_icb_cmd_valid_404;
  wire     tmp_icb_cmd_ready_404;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_404 (
    .i_vld(tmp_icb_cmd_valid_403), 
    .i_rdy(tmp_icb_cmd_ready_403), 
    .i_dat(tmp_icb_cmd_pack_403),
    .o_vld(tmp_icb_cmd_valid_404), 
    .o_rdy(delay_stage_select[404] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_404), 
    .o_dat(tmp_icb_cmd_pack_404),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_405;
  wire     tmp_icb_cmd_valid_405;
  wire     tmp_icb_cmd_ready_405;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_405 (
    .i_vld(tmp_icb_cmd_valid_404), 
    .i_rdy(tmp_icb_cmd_ready_404), 
    .i_dat(tmp_icb_cmd_pack_404),
    .o_vld(tmp_icb_cmd_valid_405), 
    .o_rdy(delay_stage_select[405] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_405), 
    .o_dat(tmp_icb_cmd_pack_405),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_406;
  wire     tmp_icb_cmd_valid_406;
  wire     tmp_icb_cmd_ready_406;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_406 (
    .i_vld(tmp_icb_cmd_valid_405), 
    .i_rdy(tmp_icb_cmd_ready_405), 
    .i_dat(tmp_icb_cmd_pack_405),
    .o_vld(tmp_icb_cmd_valid_406), 
    .o_rdy(delay_stage_select[406] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_406), 
    .o_dat(tmp_icb_cmd_pack_406),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_407;
  wire     tmp_icb_cmd_valid_407;
  wire     tmp_icb_cmd_ready_407;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_407 (
    .i_vld(tmp_icb_cmd_valid_406), 
    .i_rdy(tmp_icb_cmd_ready_406), 
    .i_dat(tmp_icb_cmd_pack_406),
    .o_vld(tmp_icb_cmd_valid_407), 
    .o_rdy(delay_stage_select[407] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_407), 
    .o_dat(tmp_icb_cmd_pack_407),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_408;
  wire     tmp_icb_cmd_valid_408;
  wire     tmp_icb_cmd_ready_408;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_408 (
    .i_vld(tmp_icb_cmd_valid_407), 
    .i_rdy(tmp_icb_cmd_ready_407), 
    .i_dat(tmp_icb_cmd_pack_407),
    .o_vld(tmp_icb_cmd_valid_408), 
    .o_rdy(delay_stage_select[408] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_408), 
    .o_dat(tmp_icb_cmd_pack_408),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_409;
  wire     tmp_icb_cmd_valid_409;
  wire     tmp_icb_cmd_ready_409;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_409 (
    .i_vld(tmp_icb_cmd_valid_408), 
    .i_rdy(tmp_icb_cmd_ready_408), 
    .i_dat(tmp_icb_cmd_pack_408),
    .o_vld(tmp_icb_cmd_valid_409), 
    .o_rdy(delay_stage_select[409] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_409), 
    .o_dat(tmp_icb_cmd_pack_409),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_410;
  wire     tmp_icb_cmd_valid_410;
  wire     tmp_icb_cmd_ready_410;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_410 (
    .i_vld(tmp_icb_cmd_valid_409), 
    .i_rdy(tmp_icb_cmd_ready_409), 
    .i_dat(tmp_icb_cmd_pack_409),
    .o_vld(tmp_icb_cmd_valid_410), 
    .o_rdy(delay_stage_select[410] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_410), 
    .o_dat(tmp_icb_cmd_pack_410),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_411;
  wire     tmp_icb_cmd_valid_411;
  wire     tmp_icb_cmd_ready_411;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_411 (
    .i_vld(tmp_icb_cmd_valid_410), 
    .i_rdy(tmp_icb_cmd_ready_410), 
    .i_dat(tmp_icb_cmd_pack_410),
    .o_vld(tmp_icb_cmd_valid_411), 
    .o_rdy(delay_stage_select[411] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_411), 
    .o_dat(tmp_icb_cmd_pack_411),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_412;
  wire     tmp_icb_cmd_valid_412;
  wire     tmp_icb_cmd_ready_412;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_412 (
    .i_vld(tmp_icb_cmd_valid_411), 
    .i_rdy(tmp_icb_cmd_ready_411), 
    .i_dat(tmp_icb_cmd_pack_411),
    .o_vld(tmp_icb_cmd_valid_412), 
    .o_rdy(delay_stage_select[412] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_412), 
    .o_dat(tmp_icb_cmd_pack_412),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_413;
  wire     tmp_icb_cmd_valid_413;
  wire     tmp_icb_cmd_ready_413;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_413 (
    .i_vld(tmp_icb_cmd_valid_412), 
    .i_rdy(tmp_icb_cmd_ready_412), 
    .i_dat(tmp_icb_cmd_pack_412),
    .o_vld(tmp_icb_cmd_valid_413), 
    .o_rdy(delay_stage_select[413] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_413), 
    .o_dat(tmp_icb_cmd_pack_413),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_414;
  wire     tmp_icb_cmd_valid_414;
  wire     tmp_icb_cmd_ready_414;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_414 (
    .i_vld(tmp_icb_cmd_valid_413), 
    .i_rdy(tmp_icb_cmd_ready_413), 
    .i_dat(tmp_icb_cmd_pack_413),
    .o_vld(tmp_icb_cmd_valid_414), 
    .o_rdy(delay_stage_select[414] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_414), 
    .o_dat(tmp_icb_cmd_pack_414),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_415;
  wire     tmp_icb_cmd_valid_415;
  wire     tmp_icb_cmd_ready_415;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_415 (
    .i_vld(tmp_icb_cmd_valid_414), 
    .i_rdy(tmp_icb_cmd_ready_414), 
    .i_dat(tmp_icb_cmd_pack_414),
    .o_vld(tmp_icb_cmd_valid_415), 
    .o_rdy(delay_stage_select[415] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_415), 
    .o_dat(tmp_icb_cmd_pack_415),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_416;
  wire     tmp_icb_cmd_valid_416;
  wire     tmp_icb_cmd_ready_416;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_416 (
    .i_vld(tmp_icb_cmd_valid_415), 
    .i_rdy(tmp_icb_cmd_ready_415), 
    .i_dat(tmp_icb_cmd_pack_415),
    .o_vld(tmp_icb_cmd_valid_416), 
    .o_rdy(delay_stage_select[416] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_416), 
    .o_dat(tmp_icb_cmd_pack_416),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_417;
  wire     tmp_icb_cmd_valid_417;
  wire     tmp_icb_cmd_ready_417;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_417 (
    .i_vld(tmp_icb_cmd_valid_416), 
    .i_rdy(tmp_icb_cmd_ready_416), 
    .i_dat(tmp_icb_cmd_pack_416),
    .o_vld(tmp_icb_cmd_valid_417), 
    .o_rdy(delay_stage_select[417] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_417), 
    .o_dat(tmp_icb_cmd_pack_417),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_418;
  wire     tmp_icb_cmd_valid_418;
  wire     tmp_icb_cmd_ready_418;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_418 (
    .i_vld(tmp_icb_cmd_valid_417), 
    .i_rdy(tmp_icb_cmd_ready_417), 
    .i_dat(tmp_icb_cmd_pack_417),
    .o_vld(tmp_icb_cmd_valid_418), 
    .o_rdy(delay_stage_select[418] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_418), 
    .o_dat(tmp_icb_cmd_pack_418),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_419;
  wire     tmp_icb_cmd_valid_419;
  wire     tmp_icb_cmd_ready_419;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_419 (
    .i_vld(tmp_icb_cmd_valid_418), 
    .i_rdy(tmp_icb_cmd_ready_418), 
    .i_dat(tmp_icb_cmd_pack_418),
    .o_vld(tmp_icb_cmd_valid_419), 
    .o_rdy(delay_stage_select[419] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_419), 
    .o_dat(tmp_icb_cmd_pack_419),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_420;
  wire     tmp_icb_cmd_valid_420;
  wire     tmp_icb_cmd_ready_420;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_420 (
    .i_vld(tmp_icb_cmd_valid_419), 
    .i_rdy(tmp_icb_cmd_ready_419), 
    .i_dat(tmp_icb_cmd_pack_419),
    .o_vld(tmp_icb_cmd_valid_420), 
    .o_rdy(delay_stage_select[420] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_420), 
    .o_dat(tmp_icb_cmd_pack_420),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_421;
  wire     tmp_icb_cmd_valid_421;
  wire     tmp_icb_cmd_ready_421;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_421 (
    .i_vld(tmp_icb_cmd_valid_420), 
    .i_rdy(tmp_icb_cmd_ready_420), 
    .i_dat(tmp_icb_cmd_pack_420),
    .o_vld(tmp_icb_cmd_valid_421), 
    .o_rdy(delay_stage_select[421] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_421), 
    .o_dat(tmp_icb_cmd_pack_421),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_422;
  wire     tmp_icb_cmd_valid_422;
  wire     tmp_icb_cmd_ready_422;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_422 (
    .i_vld(tmp_icb_cmd_valid_421), 
    .i_rdy(tmp_icb_cmd_ready_421), 
    .i_dat(tmp_icb_cmd_pack_421),
    .o_vld(tmp_icb_cmd_valid_422), 
    .o_rdy(delay_stage_select[422] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_422), 
    .o_dat(tmp_icb_cmd_pack_422),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_423;
  wire     tmp_icb_cmd_valid_423;
  wire     tmp_icb_cmd_ready_423;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_423 (
    .i_vld(tmp_icb_cmd_valid_422), 
    .i_rdy(tmp_icb_cmd_ready_422), 
    .i_dat(tmp_icb_cmd_pack_422),
    .o_vld(tmp_icb_cmd_valid_423), 
    .o_rdy(delay_stage_select[423] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_423), 
    .o_dat(tmp_icb_cmd_pack_423),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_424;
  wire     tmp_icb_cmd_valid_424;
  wire     tmp_icb_cmd_ready_424;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_424 (
    .i_vld(tmp_icb_cmd_valid_423), 
    .i_rdy(tmp_icb_cmd_ready_423), 
    .i_dat(tmp_icb_cmd_pack_423),
    .o_vld(tmp_icb_cmd_valid_424), 
    .o_rdy(delay_stage_select[424] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_424), 
    .o_dat(tmp_icb_cmd_pack_424),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_425;
  wire     tmp_icb_cmd_valid_425;
  wire     tmp_icb_cmd_ready_425;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_425 (
    .i_vld(tmp_icb_cmd_valid_424), 
    .i_rdy(tmp_icb_cmd_ready_424), 
    .i_dat(tmp_icb_cmd_pack_424),
    .o_vld(tmp_icb_cmd_valid_425), 
    .o_rdy(delay_stage_select[425] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_425), 
    .o_dat(tmp_icb_cmd_pack_425),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_426;
  wire     tmp_icb_cmd_valid_426;
  wire     tmp_icb_cmd_ready_426;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_426 (
    .i_vld(tmp_icb_cmd_valid_425), 
    .i_rdy(tmp_icb_cmd_ready_425), 
    .i_dat(tmp_icb_cmd_pack_425),
    .o_vld(tmp_icb_cmd_valid_426), 
    .o_rdy(delay_stage_select[426] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_426), 
    .o_dat(tmp_icb_cmd_pack_426),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_427;
  wire     tmp_icb_cmd_valid_427;
  wire     tmp_icb_cmd_ready_427;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_427 (
    .i_vld(tmp_icb_cmd_valid_426), 
    .i_rdy(tmp_icb_cmd_ready_426), 
    .i_dat(tmp_icb_cmd_pack_426),
    .o_vld(tmp_icb_cmd_valid_427), 
    .o_rdy(delay_stage_select[427] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_427), 
    .o_dat(tmp_icb_cmd_pack_427),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_428;
  wire     tmp_icb_cmd_valid_428;
  wire     tmp_icb_cmd_ready_428;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_428 (
    .i_vld(tmp_icb_cmd_valid_427), 
    .i_rdy(tmp_icb_cmd_ready_427), 
    .i_dat(tmp_icb_cmd_pack_427),
    .o_vld(tmp_icb_cmd_valid_428), 
    .o_rdy(delay_stage_select[428] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_428), 
    .o_dat(tmp_icb_cmd_pack_428),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_429;
  wire     tmp_icb_cmd_valid_429;
  wire     tmp_icb_cmd_ready_429;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_429 (
    .i_vld(tmp_icb_cmd_valid_428), 
    .i_rdy(tmp_icb_cmd_ready_428), 
    .i_dat(tmp_icb_cmd_pack_428),
    .o_vld(tmp_icb_cmd_valid_429), 
    .o_rdy(delay_stage_select[429] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_429), 
    .o_dat(tmp_icb_cmd_pack_429),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_430;
  wire     tmp_icb_cmd_valid_430;
  wire     tmp_icb_cmd_ready_430;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_430 (
    .i_vld(tmp_icb_cmd_valid_429), 
    .i_rdy(tmp_icb_cmd_ready_429), 
    .i_dat(tmp_icb_cmd_pack_429),
    .o_vld(tmp_icb_cmd_valid_430), 
    .o_rdy(delay_stage_select[430] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_430), 
    .o_dat(tmp_icb_cmd_pack_430),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_431;
  wire     tmp_icb_cmd_valid_431;
  wire     tmp_icb_cmd_ready_431;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_431 (
    .i_vld(tmp_icb_cmd_valid_430), 
    .i_rdy(tmp_icb_cmd_ready_430), 
    .i_dat(tmp_icb_cmd_pack_430),
    .o_vld(tmp_icb_cmd_valid_431), 
    .o_rdy(delay_stage_select[431] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_431), 
    .o_dat(tmp_icb_cmd_pack_431),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_432;
  wire     tmp_icb_cmd_valid_432;
  wire     tmp_icb_cmd_ready_432;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_432 (
    .i_vld(tmp_icb_cmd_valid_431), 
    .i_rdy(tmp_icb_cmd_ready_431), 
    .i_dat(tmp_icb_cmd_pack_431),
    .o_vld(tmp_icb_cmd_valid_432), 
    .o_rdy(delay_stage_select[432] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_432), 
    .o_dat(tmp_icb_cmd_pack_432),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_433;
  wire     tmp_icb_cmd_valid_433;
  wire     tmp_icb_cmd_ready_433;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_433 (
    .i_vld(tmp_icb_cmd_valid_432), 
    .i_rdy(tmp_icb_cmd_ready_432), 
    .i_dat(tmp_icb_cmd_pack_432),
    .o_vld(tmp_icb_cmd_valid_433), 
    .o_rdy(delay_stage_select[433] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_433), 
    .o_dat(tmp_icb_cmd_pack_433),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_434;
  wire     tmp_icb_cmd_valid_434;
  wire     tmp_icb_cmd_ready_434;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_434 (
    .i_vld(tmp_icb_cmd_valid_433), 
    .i_rdy(tmp_icb_cmd_ready_433), 
    .i_dat(tmp_icb_cmd_pack_433),
    .o_vld(tmp_icb_cmd_valid_434), 
    .o_rdy(delay_stage_select[434] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_434), 
    .o_dat(tmp_icb_cmd_pack_434),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_435;
  wire     tmp_icb_cmd_valid_435;
  wire     tmp_icb_cmd_ready_435;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_435 (
    .i_vld(tmp_icb_cmd_valid_434), 
    .i_rdy(tmp_icb_cmd_ready_434), 
    .i_dat(tmp_icb_cmd_pack_434),
    .o_vld(tmp_icb_cmd_valid_435), 
    .o_rdy(delay_stage_select[435] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_435), 
    .o_dat(tmp_icb_cmd_pack_435),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_436;
  wire     tmp_icb_cmd_valid_436;
  wire     tmp_icb_cmd_ready_436;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_436 (
    .i_vld(tmp_icb_cmd_valid_435), 
    .i_rdy(tmp_icb_cmd_ready_435), 
    .i_dat(tmp_icb_cmd_pack_435),
    .o_vld(tmp_icb_cmd_valid_436), 
    .o_rdy(delay_stage_select[436] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_436), 
    .o_dat(tmp_icb_cmd_pack_436),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_437;
  wire     tmp_icb_cmd_valid_437;
  wire     tmp_icb_cmd_ready_437;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_437 (
    .i_vld(tmp_icb_cmd_valid_436), 
    .i_rdy(tmp_icb_cmd_ready_436), 
    .i_dat(tmp_icb_cmd_pack_436),
    .o_vld(tmp_icb_cmd_valid_437), 
    .o_rdy(delay_stage_select[437] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_437), 
    .o_dat(tmp_icb_cmd_pack_437),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_438;
  wire     tmp_icb_cmd_valid_438;
  wire     tmp_icb_cmd_ready_438;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_438 (
    .i_vld(tmp_icb_cmd_valid_437), 
    .i_rdy(tmp_icb_cmd_ready_437), 
    .i_dat(tmp_icb_cmd_pack_437),
    .o_vld(tmp_icb_cmd_valid_438), 
    .o_rdy(delay_stage_select[438] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_438), 
    .o_dat(tmp_icb_cmd_pack_438),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_439;
  wire     tmp_icb_cmd_valid_439;
  wire     tmp_icb_cmd_ready_439;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_439 (
    .i_vld(tmp_icb_cmd_valid_438), 
    .i_rdy(tmp_icb_cmd_ready_438), 
    .i_dat(tmp_icb_cmd_pack_438),
    .o_vld(tmp_icb_cmd_valid_439), 
    .o_rdy(delay_stage_select[439] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_439), 
    .o_dat(tmp_icb_cmd_pack_439),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_440;
  wire     tmp_icb_cmd_valid_440;
  wire     tmp_icb_cmd_ready_440;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_440 (
    .i_vld(tmp_icb_cmd_valid_439), 
    .i_rdy(tmp_icb_cmd_ready_439), 
    .i_dat(tmp_icb_cmd_pack_439),
    .o_vld(tmp_icb_cmd_valid_440), 
    .o_rdy(delay_stage_select[440] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_440), 
    .o_dat(tmp_icb_cmd_pack_440),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_441;
  wire     tmp_icb_cmd_valid_441;
  wire     tmp_icb_cmd_ready_441;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_441 (
    .i_vld(tmp_icb_cmd_valid_440), 
    .i_rdy(tmp_icb_cmd_ready_440), 
    .i_dat(tmp_icb_cmd_pack_440),
    .o_vld(tmp_icb_cmd_valid_441), 
    .o_rdy(delay_stage_select[441] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_441), 
    .o_dat(tmp_icb_cmd_pack_441),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_442;
  wire     tmp_icb_cmd_valid_442;
  wire     tmp_icb_cmd_ready_442;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_442 (
    .i_vld(tmp_icb_cmd_valid_441), 
    .i_rdy(tmp_icb_cmd_ready_441), 
    .i_dat(tmp_icb_cmd_pack_441),
    .o_vld(tmp_icb_cmd_valid_442), 
    .o_rdy(delay_stage_select[442] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_442), 
    .o_dat(tmp_icb_cmd_pack_442),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_443;
  wire     tmp_icb_cmd_valid_443;
  wire     tmp_icb_cmd_ready_443;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_443 (
    .i_vld(tmp_icb_cmd_valid_442), 
    .i_rdy(tmp_icb_cmd_ready_442), 
    .i_dat(tmp_icb_cmd_pack_442),
    .o_vld(tmp_icb_cmd_valid_443), 
    .o_rdy(delay_stage_select[443] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_443), 
    .o_dat(tmp_icb_cmd_pack_443),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_444;
  wire     tmp_icb_cmd_valid_444;
  wire     tmp_icb_cmd_ready_444;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_444 (
    .i_vld(tmp_icb_cmd_valid_443), 
    .i_rdy(tmp_icb_cmd_ready_443), 
    .i_dat(tmp_icb_cmd_pack_443),
    .o_vld(tmp_icb_cmd_valid_444), 
    .o_rdy(delay_stage_select[444] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_444), 
    .o_dat(tmp_icb_cmd_pack_444),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_445;
  wire     tmp_icb_cmd_valid_445;
  wire     tmp_icb_cmd_ready_445;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_445 (
    .i_vld(tmp_icb_cmd_valid_444), 
    .i_rdy(tmp_icb_cmd_ready_444), 
    .i_dat(tmp_icb_cmd_pack_444),
    .o_vld(tmp_icb_cmd_valid_445), 
    .o_rdy(delay_stage_select[445] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_445), 
    .o_dat(tmp_icb_cmd_pack_445),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_446;
  wire     tmp_icb_cmd_valid_446;
  wire     tmp_icb_cmd_ready_446;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_446 (
    .i_vld(tmp_icb_cmd_valid_445), 
    .i_rdy(tmp_icb_cmd_ready_445), 
    .i_dat(tmp_icb_cmd_pack_445),
    .o_vld(tmp_icb_cmd_valid_446), 
    .o_rdy(delay_stage_select[446] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_446), 
    .o_dat(tmp_icb_cmd_pack_446),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_447;
  wire     tmp_icb_cmd_valid_447;
  wire     tmp_icb_cmd_ready_447;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_447 (
    .i_vld(tmp_icb_cmd_valid_446), 
    .i_rdy(tmp_icb_cmd_ready_446), 
    .i_dat(tmp_icb_cmd_pack_446),
    .o_vld(tmp_icb_cmd_valid_447), 
    .o_rdy(delay_stage_select[447] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_447), 
    .o_dat(tmp_icb_cmd_pack_447),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_448;
  wire     tmp_icb_cmd_valid_448;
  wire     tmp_icb_cmd_ready_448;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_448 (
    .i_vld(tmp_icb_cmd_valid_447), 
    .i_rdy(tmp_icb_cmd_ready_447), 
    .i_dat(tmp_icb_cmd_pack_447),
    .o_vld(tmp_icb_cmd_valid_448), 
    .o_rdy(delay_stage_select[448] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_448), 
    .o_dat(tmp_icb_cmd_pack_448),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_449;
  wire     tmp_icb_cmd_valid_449;
  wire     tmp_icb_cmd_ready_449;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_449 (
    .i_vld(tmp_icb_cmd_valid_448), 
    .i_rdy(tmp_icb_cmd_ready_448), 
    .i_dat(tmp_icb_cmd_pack_448),
    .o_vld(tmp_icb_cmd_valid_449), 
    .o_rdy(delay_stage_select[449] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_449), 
    .o_dat(tmp_icb_cmd_pack_449),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_450;
  wire     tmp_icb_cmd_valid_450;
  wire     tmp_icb_cmd_ready_450;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_450 (
    .i_vld(tmp_icb_cmd_valid_449), 
    .i_rdy(tmp_icb_cmd_ready_449), 
    .i_dat(tmp_icb_cmd_pack_449),
    .o_vld(tmp_icb_cmd_valid_450), 
    .o_rdy(delay_stage_select[450] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_450), 
    .o_dat(tmp_icb_cmd_pack_450),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_451;
  wire     tmp_icb_cmd_valid_451;
  wire     tmp_icb_cmd_ready_451;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_451 (
    .i_vld(tmp_icb_cmd_valid_450), 
    .i_rdy(tmp_icb_cmd_ready_450), 
    .i_dat(tmp_icb_cmd_pack_450),
    .o_vld(tmp_icb_cmd_valid_451), 
    .o_rdy(delay_stage_select[451] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_451), 
    .o_dat(tmp_icb_cmd_pack_451),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_452;
  wire     tmp_icb_cmd_valid_452;
  wire     tmp_icb_cmd_ready_452;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_452 (
    .i_vld(tmp_icb_cmd_valid_451), 
    .i_rdy(tmp_icb_cmd_ready_451), 
    .i_dat(tmp_icb_cmd_pack_451),
    .o_vld(tmp_icb_cmd_valid_452), 
    .o_rdy(delay_stage_select[452] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_452), 
    .o_dat(tmp_icb_cmd_pack_452),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_453;
  wire     tmp_icb_cmd_valid_453;
  wire     tmp_icb_cmd_ready_453;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_453 (
    .i_vld(tmp_icb_cmd_valid_452), 
    .i_rdy(tmp_icb_cmd_ready_452), 
    .i_dat(tmp_icb_cmd_pack_452),
    .o_vld(tmp_icb_cmd_valid_453), 
    .o_rdy(delay_stage_select[453] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_453), 
    .o_dat(tmp_icb_cmd_pack_453),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_454;
  wire     tmp_icb_cmd_valid_454;
  wire     tmp_icb_cmd_ready_454;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_454 (
    .i_vld(tmp_icb_cmd_valid_453), 
    .i_rdy(tmp_icb_cmd_ready_453), 
    .i_dat(tmp_icb_cmd_pack_453),
    .o_vld(tmp_icb_cmd_valid_454), 
    .o_rdy(delay_stage_select[454] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_454), 
    .o_dat(tmp_icb_cmd_pack_454),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_455;
  wire     tmp_icb_cmd_valid_455;
  wire     tmp_icb_cmd_ready_455;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_455 (
    .i_vld(tmp_icb_cmd_valid_454), 
    .i_rdy(tmp_icb_cmd_ready_454), 
    .i_dat(tmp_icb_cmd_pack_454),
    .o_vld(tmp_icb_cmd_valid_455), 
    .o_rdy(delay_stage_select[455] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_455), 
    .o_dat(tmp_icb_cmd_pack_455),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_456;
  wire     tmp_icb_cmd_valid_456;
  wire     tmp_icb_cmd_ready_456;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_456 (
    .i_vld(tmp_icb_cmd_valid_455), 
    .i_rdy(tmp_icb_cmd_ready_455), 
    .i_dat(tmp_icb_cmd_pack_455),
    .o_vld(tmp_icb_cmd_valid_456), 
    .o_rdy(delay_stage_select[456] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_456), 
    .o_dat(tmp_icb_cmd_pack_456),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_457;
  wire     tmp_icb_cmd_valid_457;
  wire     tmp_icb_cmd_ready_457;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_457 (
    .i_vld(tmp_icb_cmd_valid_456), 
    .i_rdy(tmp_icb_cmd_ready_456), 
    .i_dat(tmp_icb_cmd_pack_456),
    .o_vld(tmp_icb_cmd_valid_457), 
    .o_rdy(delay_stage_select[457] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_457), 
    .o_dat(tmp_icb_cmd_pack_457),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_458;
  wire     tmp_icb_cmd_valid_458;
  wire     tmp_icb_cmd_ready_458;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_458 (
    .i_vld(tmp_icb_cmd_valid_457), 
    .i_rdy(tmp_icb_cmd_ready_457), 
    .i_dat(tmp_icb_cmd_pack_457),
    .o_vld(tmp_icb_cmd_valid_458), 
    .o_rdy(delay_stage_select[458] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_458), 
    .o_dat(tmp_icb_cmd_pack_458),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_459;
  wire     tmp_icb_cmd_valid_459;
  wire     tmp_icb_cmd_ready_459;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_459 (
    .i_vld(tmp_icb_cmd_valid_458), 
    .i_rdy(tmp_icb_cmd_ready_458), 
    .i_dat(tmp_icb_cmd_pack_458),
    .o_vld(tmp_icb_cmd_valid_459), 
    .o_rdy(delay_stage_select[459] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_459), 
    .o_dat(tmp_icb_cmd_pack_459),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_460;
  wire     tmp_icb_cmd_valid_460;
  wire     tmp_icb_cmd_ready_460;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_460 (
    .i_vld(tmp_icb_cmd_valid_459), 
    .i_rdy(tmp_icb_cmd_ready_459), 
    .i_dat(tmp_icb_cmd_pack_459),
    .o_vld(tmp_icb_cmd_valid_460), 
    .o_rdy(delay_stage_select[460] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_460), 
    .o_dat(tmp_icb_cmd_pack_460),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_461;
  wire     tmp_icb_cmd_valid_461;
  wire     tmp_icb_cmd_ready_461;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_461 (
    .i_vld(tmp_icb_cmd_valid_460), 
    .i_rdy(tmp_icb_cmd_ready_460), 
    .i_dat(tmp_icb_cmd_pack_460),
    .o_vld(tmp_icb_cmd_valid_461), 
    .o_rdy(delay_stage_select[461] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_461), 
    .o_dat(tmp_icb_cmd_pack_461),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_462;
  wire     tmp_icb_cmd_valid_462;
  wire     tmp_icb_cmd_ready_462;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_462 (
    .i_vld(tmp_icb_cmd_valid_461), 
    .i_rdy(tmp_icb_cmd_ready_461), 
    .i_dat(tmp_icb_cmd_pack_461),
    .o_vld(tmp_icb_cmd_valid_462), 
    .o_rdy(delay_stage_select[462] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_462), 
    .o_dat(tmp_icb_cmd_pack_462),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_463;
  wire     tmp_icb_cmd_valid_463;
  wire     tmp_icb_cmd_ready_463;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_463 (
    .i_vld(tmp_icb_cmd_valid_462), 
    .i_rdy(tmp_icb_cmd_ready_462), 
    .i_dat(tmp_icb_cmd_pack_462),
    .o_vld(tmp_icb_cmd_valid_463), 
    .o_rdy(delay_stage_select[463] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_463), 
    .o_dat(tmp_icb_cmd_pack_463),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_464;
  wire     tmp_icb_cmd_valid_464;
  wire     tmp_icb_cmd_ready_464;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_464 (
    .i_vld(tmp_icb_cmd_valid_463), 
    .i_rdy(tmp_icb_cmd_ready_463), 
    .i_dat(tmp_icb_cmd_pack_463),
    .o_vld(tmp_icb_cmd_valid_464), 
    .o_rdy(delay_stage_select[464] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_464), 
    .o_dat(tmp_icb_cmd_pack_464),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_465;
  wire     tmp_icb_cmd_valid_465;
  wire     tmp_icb_cmd_ready_465;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_465 (
    .i_vld(tmp_icb_cmd_valid_464), 
    .i_rdy(tmp_icb_cmd_ready_464), 
    .i_dat(tmp_icb_cmd_pack_464),
    .o_vld(tmp_icb_cmd_valid_465), 
    .o_rdy(delay_stage_select[465] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_465), 
    .o_dat(tmp_icb_cmd_pack_465),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_466;
  wire     tmp_icb_cmd_valid_466;
  wire     tmp_icb_cmd_ready_466;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_466 (
    .i_vld(tmp_icb_cmd_valid_465), 
    .i_rdy(tmp_icb_cmd_ready_465), 
    .i_dat(tmp_icb_cmd_pack_465),
    .o_vld(tmp_icb_cmd_valid_466), 
    .o_rdy(delay_stage_select[466] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_466), 
    .o_dat(tmp_icb_cmd_pack_466),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_467;
  wire     tmp_icb_cmd_valid_467;
  wire     tmp_icb_cmd_ready_467;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_467 (
    .i_vld(tmp_icb_cmd_valid_466), 
    .i_rdy(tmp_icb_cmd_ready_466), 
    .i_dat(tmp_icb_cmd_pack_466),
    .o_vld(tmp_icb_cmd_valid_467), 
    .o_rdy(delay_stage_select[467] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_467), 
    .o_dat(tmp_icb_cmd_pack_467),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_468;
  wire     tmp_icb_cmd_valid_468;
  wire     tmp_icb_cmd_ready_468;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_468 (
    .i_vld(tmp_icb_cmd_valid_467), 
    .i_rdy(tmp_icb_cmd_ready_467), 
    .i_dat(tmp_icb_cmd_pack_467),
    .o_vld(tmp_icb_cmd_valid_468), 
    .o_rdy(delay_stage_select[468] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_468), 
    .o_dat(tmp_icb_cmd_pack_468),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_469;
  wire     tmp_icb_cmd_valid_469;
  wire     tmp_icb_cmd_ready_469;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_469 (
    .i_vld(tmp_icb_cmd_valid_468), 
    .i_rdy(tmp_icb_cmd_ready_468), 
    .i_dat(tmp_icb_cmd_pack_468),
    .o_vld(tmp_icb_cmd_valid_469), 
    .o_rdy(delay_stage_select[469] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_469), 
    .o_dat(tmp_icb_cmd_pack_469),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_470;
  wire     tmp_icb_cmd_valid_470;
  wire     tmp_icb_cmd_ready_470;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_470 (
    .i_vld(tmp_icb_cmd_valid_469), 
    .i_rdy(tmp_icb_cmd_ready_469), 
    .i_dat(tmp_icb_cmd_pack_469),
    .o_vld(tmp_icb_cmd_valid_470), 
    .o_rdy(delay_stage_select[470] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_470), 
    .o_dat(tmp_icb_cmd_pack_470),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_471;
  wire     tmp_icb_cmd_valid_471;
  wire     tmp_icb_cmd_ready_471;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_471 (
    .i_vld(tmp_icb_cmd_valid_470), 
    .i_rdy(tmp_icb_cmd_ready_470), 
    .i_dat(tmp_icb_cmd_pack_470),
    .o_vld(tmp_icb_cmd_valid_471), 
    .o_rdy(delay_stage_select[471] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_471), 
    .o_dat(tmp_icb_cmd_pack_471),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_472;
  wire     tmp_icb_cmd_valid_472;
  wire     tmp_icb_cmd_ready_472;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_472 (
    .i_vld(tmp_icb_cmd_valid_471), 
    .i_rdy(tmp_icb_cmd_ready_471), 
    .i_dat(tmp_icb_cmd_pack_471),
    .o_vld(tmp_icb_cmd_valid_472), 
    .o_rdy(delay_stage_select[472] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_472), 
    .o_dat(tmp_icb_cmd_pack_472),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_473;
  wire     tmp_icb_cmd_valid_473;
  wire     tmp_icb_cmd_ready_473;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_473 (
    .i_vld(tmp_icb_cmd_valid_472), 
    .i_rdy(tmp_icb_cmd_ready_472), 
    .i_dat(tmp_icb_cmd_pack_472),
    .o_vld(tmp_icb_cmd_valid_473), 
    .o_rdy(delay_stage_select[473] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_473), 
    .o_dat(tmp_icb_cmd_pack_473),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_474;
  wire     tmp_icb_cmd_valid_474;
  wire     tmp_icb_cmd_ready_474;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_474 (
    .i_vld(tmp_icb_cmd_valid_473), 
    .i_rdy(tmp_icb_cmd_ready_473), 
    .i_dat(tmp_icb_cmd_pack_473),
    .o_vld(tmp_icb_cmd_valid_474), 
    .o_rdy(delay_stage_select[474] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_474), 
    .o_dat(tmp_icb_cmd_pack_474),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_475;
  wire     tmp_icb_cmd_valid_475;
  wire     tmp_icb_cmd_ready_475;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_475 (
    .i_vld(tmp_icb_cmd_valid_474), 
    .i_rdy(tmp_icb_cmd_ready_474), 
    .i_dat(tmp_icb_cmd_pack_474),
    .o_vld(tmp_icb_cmd_valid_475), 
    .o_rdy(delay_stage_select[475] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_475), 
    .o_dat(tmp_icb_cmd_pack_475),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_476;
  wire     tmp_icb_cmd_valid_476;
  wire     tmp_icb_cmd_ready_476;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_476 (
    .i_vld(tmp_icb_cmd_valid_475), 
    .i_rdy(tmp_icb_cmd_ready_475), 
    .i_dat(tmp_icb_cmd_pack_475),
    .o_vld(tmp_icb_cmd_valid_476), 
    .o_rdy(delay_stage_select[476] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_476), 
    .o_dat(tmp_icb_cmd_pack_476),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_477;
  wire     tmp_icb_cmd_valid_477;
  wire     tmp_icb_cmd_ready_477;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_477 (
    .i_vld(tmp_icb_cmd_valid_476), 
    .i_rdy(tmp_icb_cmd_ready_476), 
    .i_dat(tmp_icb_cmd_pack_476),
    .o_vld(tmp_icb_cmd_valid_477), 
    .o_rdy(delay_stage_select[477] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_477), 
    .o_dat(tmp_icb_cmd_pack_477),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_478;
  wire     tmp_icb_cmd_valid_478;
  wire     tmp_icb_cmd_ready_478;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_478 (
    .i_vld(tmp_icb_cmd_valid_477), 
    .i_rdy(tmp_icb_cmd_ready_477), 
    .i_dat(tmp_icb_cmd_pack_477),
    .o_vld(tmp_icb_cmd_valid_478), 
    .o_rdy(delay_stage_select[478] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_478), 
    .o_dat(tmp_icb_cmd_pack_478),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_479;
  wire     tmp_icb_cmd_valid_479;
  wire     tmp_icb_cmd_ready_479;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_479 (
    .i_vld(tmp_icb_cmd_valid_478), 
    .i_rdy(tmp_icb_cmd_ready_478), 
    .i_dat(tmp_icb_cmd_pack_478),
    .o_vld(tmp_icb_cmd_valid_479), 
    .o_rdy(delay_stage_select[479] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_479), 
    .o_dat(tmp_icb_cmd_pack_479),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_480;
  wire     tmp_icb_cmd_valid_480;
  wire     tmp_icb_cmd_ready_480;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_480 (
    .i_vld(tmp_icb_cmd_valid_479), 
    .i_rdy(tmp_icb_cmd_ready_479), 
    .i_dat(tmp_icb_cmd_pack_479),
    .o_vld(tmp_icb_cmd_valid_480), 
    .o_rdy(delay_stage_select[480] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_480), 
    .o_dat(tmp_icb_cmd_pack_480),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_481;
  wire     tmp_icb_cmd_valid_481;
  wire     tmp_icb_cmd_ready_481;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_481 (
    .i_vld(tmp_icb_cmd_valid_480), 
    .i_rdy(tmp_icb_cmd_ready_480), 
    .i_dat(tmp_icb_cmd_pack_480),
    .o_vld(tmp_icb_cmd_valid_481), 
    .o_rdy(delay_stage_select[481] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_481), 
    .o_dat(tmp_icb_cmd_pack_481),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_482;
  wire     tmp_icb_cmd_valid_482;
  wire     tmp_icb_cmd_ready_482;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_482 (
    .i_vld(tmp_icb_cmd_valid_481), 
    .i_rdy(tmp_icb_cmd_ready_481), 
    .i_dat(tmp_icb_cmd_pack_481),
    .o_vld(tmp_icb_cmd_valid_482), 
    .o_rdy(delay_stage_select[482] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_482), 
    .o_dat(tmp_icb_cmd_pack_482),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_483;
  wire     tmp_icb_cmd_valid_483;
  wire     tmp_icb_cmd_ready_483;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_483 (
    .i_vld(tmp_icb_cmd_valid_482), 
    .i_rdy(tmp_icb_cmd_ready_482), 
    .i_dat(tmp_icb_cmd_pack_482),
    .o_vld(tmp_icb_cmd_valid_483), 
    .o_rdy(delay_stage_select[483] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_483), 
    .o_dat(tmp_icb_cmd_pack_483),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_484;
  wire     tmp_icb_cmd_valid_484;
  wire     tmp_icb_cmd_ready_484;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_484 (
    .i_vld(tmp_icb_cmd_valid_483), 
    .i_rdy(tmp_icb_cmd_ready_483), 
    .i_dat(tmp_icb_cmd_pack_483),
    .o_vld(tmp_icb_cmd_valid_484), 
    .o_rdy(delay_stage_select[484] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_484), 
    .o_dat(tmp_icb_cmd_pack_484),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_485;
  wire     tmp_icb_cmd_valid_485;
  wire     tmp_icb_cmd_ready_485;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_485 (
    .i_vld(tmp_icb_cmd_valid_484), 
    .i_rdy(tmp_icb_cmd_ready_484), 
    .i_dat(tmp_icb_cmd_pack_484),
    .o_vld(tmp_icb_cmd_valid_485), 
    .o_rdy(delay_stage_select[485] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_485), 
    .o_dat(tmp_icb_cmd_pack_485),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_486;
  wire     tmp_icb_cmd_valid_486;
  wire     tmp_icb_cmd_ready_486;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_486 (
    .i_vld(tmp_icb_cmd_valid_485), 
    .i_rdy(tmp_icb_cmd_ready_485), 
    .i_dat(tmp_icb_cmd_pack_485),
    .o_vld(tmp_icb_cmd_valid_486), 
    .o_rdy(delay_stage_select[486] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_486), 
    .o_dat(tmp_icb_cmd_pack_486),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_487;
  wire     tmp_icb_cmd_valid_487;
  wire     tmp_icb_cmd_ready_487;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_487 (
    .i_vld(tmp_icb_cmd_valid_486), 
    .i_rdy(tmp_icb_cmd_ready_486), 
    .i_dat(tmp_icb_cmd_pack_486),
    .o_vld(tmp_icb_cmd_valid_487), 
    .o_rdy(delay_stage_select[487] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_487), 
    .o_dat(tmp_icb_cmd_pack_487),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_488;
  wire     tmp_icb_cmd_valid_488;
  wire     tmp_icb_cmd_ready_488;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_488 (
    .i_vld(tmp_icb_cmd_valid_487), 
    .i_rdy(tmp_icb_cmd_ready_487), 
    .i_dat(tmp_icb_cmd_pack_487),
    .o_vld(tmp_icb_cmd_valid_488), 
    .o_rdy(delay_stage_select[488] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_488), 
    .o_dat(tmp_icb_cmd_pack_488),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_489;
  wire     tmp_icb_cmd_valid_489;
  wire     tmp_icb_cmd_ready_489;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_489 (
    .i_vld(tmp_icb_cmd_valid_488), 
    .i_rdy(tmp_icb_cmd_ready_488), 
    .i_dat(tmp_icb_cmd_pack_488),
    .o_vld(tmp_icb_cmd_valid_489), 
    .o_rdy(delay_stage_select[489] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_489), 
    .o_dat(tmp_icb_cmd_pack_489),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_490;
  wire     tmp_icb_cmd_valid_490;
  wire     tmp_icb_cmd_ready_490;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_490 (
    .i_vld(tmp_icb_cmd_valid_489), 
    .i_rdy(tmp_icb_cmd_ready_489), 
    .i_dat(tmp_icb_cmd_pack_489),
    .o_vld(tmp_icb_cmd_valid_490), 
    .o_rdy(delay_stage_select[490] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_490), 
    .o_dat(tmp_icb_cmd_pack_490),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_491;
  wire     tmp_icb_cmd_valid_491;
  wire     tmp_icb_cmd_ready_491;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_491 (
    .i_vld(tmp_icb_cmd_valid_490), 
    .i_rdy(tmp_icb_cmd_ready_490), 
    .i_dat(tmp_icb_cmd_pack_490),
    .o_vld(tmp_icb_cmd_valid_491), 
    .o_rdy(delay_stage_select[491] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_491), 
    .o_dat(tmp_icb_cmd_pack_491),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_492;
  wire     tmp_icb_cmd_valid_492;
  wire     tmp_icb_cmd_ready_492;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_492 (
    .i_vld(tmp_icb_cmd_valid_491), 
    .i_rdy(tmp_icb_cmd_ready_491), 
    .i_dat(tmp_icb_cmd_pack_491),
    .o_vld(tmp_icb_cmd_valid_492), 
    .o_rdy(delay_stage_select[492] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_492), 
    .o_dat(tmp_icb_cmd_pack_492),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_493;
  wire     tmp_icb_cmd_valid_493;
  wire     tmp_icb_cmd_ready_493;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_493 (
    .i_vld(tmp_icb_cmd_valid_492), 
    .i_rdy(tmp_icb_cmd_ready_492), 
    .i_dat(tmp_icb_cmd_pack_492),
    .o_vld(tmp_icb_cmd_valid_493), 
    .o_rdy(delay_stage_select[493] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_493), 
    .o_dat(tmp_icb_cmd_pack_493),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_494;
  wire     tmp_icb_cmd_valid_494;
  wire     tmp_icb_cmd_ready_494;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_494 (
    .i_vld(tmp_icb_cmd_valid_493), 
    .i_rdy(tmp_icb_cmd_ready_493), 
    .i_dat(tmp_icb_cmd_pack_493),
    .o_vld(tmp_icb_cmd_valid_494), 
    .o_rdy(delay_stage_select[494] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_494), 
    .o_dat(tmp_icb_cmd_pack_494),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_495;
  wire     tmp_icb_cmd_valid_495;
  wire     tmp_icb_cmd_ready_495;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_495 (
    .i_vld(tmp_icb_cmd_valid_494), 
    .i_rdy(tmp_icb_cmd_ready_494), 
    .i_dat(tmp_icb_cmd_pack_494),
    .o_vld(tmp_icb_cmd_valid_495), 
    .o_rdy(delay_stage_select[495] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_495), 
    .o_dat(tmp_icb_cmd_pack_495),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_496;
  wire     tmp_icb_cmd_valid_496;
  wire     tmp_icb_cmd_ready_496;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_496 (
    .i_vld(tmp_icb_cmd_valid_495), 
    .i_rdy(tmp_icb_cmd_ready_495), 
    .i_dat(tmp_icb_cmd_pack_495),
    .o_vld(tmp_icb_cmd_valid_496), 
    .o_rdy(delay_stage_select[496] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_496), 
    .o_dat(tmp_icb_cmd_pack_496),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_497;
  wire     tmp_icb_cmd_valid_497;
  wire     tmp_icb_cmd_ready_497;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_497 (
    .i_vld(tmp_icb_cmd_valid_496), 
    .i_rdy(tmp_icb_cmd_ready_496), 
    .i_dat(tmp_icb_cmd_pack_496),
    .o_vld(tmp_icb_cmd_valid_497), 
    .o_rdy(delay_stage_select[497] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_497), 
    .o_dat(tmp_icb_cmd_pack_497),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_498;
  wire     tmp_icb_cmd_valid_498;
  wire     tmp_icb_cmd_ready_498;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_498 (
    .i_vld(tmp_icb_cmd_valid_497), 
    .i_rdy(tmp_icb_cmd_ready_497), 
    .i_dat(tmp_icb_cmd_pack_497),
    .o_vld(tmp_icb_cmd_valid_498), 
    .o_rdy(delay_stage_select[498] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_498), 
    .o_dat(tmp_icb_cmd_pack_498),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_499;
  wire     tmp_icb_cmd_valid_499;
  wire     tmp_icb_cmd_ready_499;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_499 (
    .i_vld(tmp_icb_cmd_valid_498), 
    .i_rdy(tmp_icb_cmd_ready_498), 
    .i_dat(tmp_icb_cmd_pack_498),
    .o_vld(tmp_icb_cmd_valid_499), 
    .o_rdy(delay_stage_select[499] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_499), 
    .o_dat(tmp_icb_cmd_pack_499),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_500;
  wire     tmp_icb_cmd_valid_500;
  wire     tmp_icb_cmd_ready_500;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_500 (
    .i_vld(tmp_icb_cmd_valid_499), 
    .i_rdy(tmp_icb_cmd_ready_499), 
    .i_dat(tmp_icb_cmd_pack_499),
    .o_vld(tmp_icb_cmd_valid_500), 
    .o_rdy(delay_stage_select[500] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_500), 
    .o_dat(tmp_icb_cmd_pack_500),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_501;
  wire     tmp_icb_cmd_valid_501;
  wire     tmp_icb_cmd_ready_501;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_501 (
    .i_vld(tmp_icb_cmd_valid_500), 
    .i_rdy(tmp_icb_cmd_ready_500), 
    .i_dat(tmp_icb_cmd_pack_500),
    .o_vld(tmp_icb_cmd_valid_501), 
    .o_rdy(delay_stage_select[501] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_501), 
    .o_dat(tmp_icb_cmd_pack_501),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_502;
  wire     tmp_icb_cmd_valid_502;
  wire     tmp_icb_cmd_ready_502;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_502 (
    .i_vld(tmp_icb_cmd_valid_501), 
    .i_rdy(tmp_icb_cmd_ready_501), 
    .i_dat(tmp_icb_cmd_pack_501),
    .o_vld(tmp_icb_cmd_valid_502), 
    .o_rdy(delay_stage_select[502] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_502), 
    .o_dat(tmp_icb_cmd_pack_502),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_503;
  wire     tmp_icb_cmd_valid_503;
  wire     tmp_icb_cmd_ready_503;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_503 (
    .i_vld(tmp_icb_cmd_valid_502), 
    .i_rdy(tmp_icb_cmd_ready_502), 
    .i_dat(tmp_icb_cmd_pack_502),
    .o_vld(tmp_icb_cmd_valid_503), 
    .o_rdy(delay_stage_select[503] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_503), 
    .o_dat(tmp_icb_cmd_pack_503),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_504;
  wire     tmp_icb_cmd_valid_504;
  wire     tmp_icb_cmd_ready_504;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_504 (
    .i_vld(tmp_icb_cmd_valid_503), 
    .i_rdy(tmp_icb_cmd_ready_503), 
    .i_dat(tmp_icb_cmd_pack_503),
    .o_vld(tmp_icb_cmd_valid_504), 
    .o_rdy(delay_stage_select[504] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_504), 
    .o_dat(tmp_icb_cmd_pack_504),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_505;
  wire     tmp_icb_cmd_valid_505;
  wire     tmp_icb_cmd_ready_505;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_505 (
    .i_vld(tmp_icb_cmd_valid_504), 
    .i_rdy(tmp_icb_cmd_ready_504), 
    .i_dat(tmp_icb_cmd_pack_504),
    .o_vld(tmp_icb_cmd_valid_505), 
    .o_rdy(delay_stage_select[505] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_505), 
    .o_dat(tmp_icb_cmd_pack_505),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_506;
  wire     tmp_icb_cmd_valid_506;
  wire     tmp_icb_cmd_ready_506;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_506 (
    .i_vld(tmp_icb_cmd_valid_505), 
    .i_rdy(tmp_icb_cmd_ready_505), 
    .i_dat(tmp_icb_cmd_pack_505),
    .o_vld(tmp_icb_cmd_valid_506), 
    .o_rdy(delay_stage_select[506] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_506), 
    .o_dat(tmp_icb_cmd_pack_506),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_507;
  wire     tmp_icb_cmd_valid_507;
  wire     tmp_icb_cmd_ready_507;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_507 (
    .i_vld(tmp_icb_cmd_valid_506), 
    .i_rdy(tmp_icb_cmd_ready_506), 
    .i_dat(tmp_icb_cmd_pack_506),
    .o_vld(tmp_icb_cmd_valid_507), 
    .o_rdy(delay_stage_select[507] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_507), 
    .o_dat(tmp_icb_cmd_pack_507),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_508;
  wire     tmp_icb_cmd_valid_508;
  wire     tmp_icb_cmd_ready_508;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_508 (
    .i_vld(tmp_icb_cmd_valid_507), 
    .i_rdy(tmp_icb_cmd_ready_507), 
    .i_dat(tmp_icb_cmd_pack_507),
    .o_vld(tmp_icb_cmd_valid_508), 
    .o_rdy(delay_stage_select[508] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_508), 
    .o_dat(tmp_icb_cmd_pack_508),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_509;
  wire     tmp_icb_cmd_valid_509;
  wire     tmp_icb_cmd_ready_509;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_509 (
    .i_vld(tmp_icb_cmd_valid_508), 
    .i_rdy(tmp_icb_cmd_ready_508), 
    .i_dat(tmp_icb_cmd_pack_508),
    .o_vld(tmp_icb_cmd_valid_509), 
    .o_rdy(delay_stage_select[509] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_509), 
    .o_dat(tmp_icb_cmd_pack_509),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_510;
  wire     tmp_icb_cmd_valid_510;
  wire     tmp_icb_cmd_ready_510;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_510 (
    .i_vld(tmp_icb_cmd_valid_509), 
    .i_rdy(tmp_icb_cmd_ready_509), 
    .i_dat(tmp_icb_cmd_pack_509),
    .o_vld(tmp_icb_cmd_valid_510), 
    .o_rdy(delay_stage_select[510] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_510), 
    .o_dat(tmp_icb_cmd_pack_510),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [BUF_CMD_PACK_W-1:0] tmp_icb_cmd_pack_511;
  wire     tmp_icb_cmd_valid_511;
  wire     tmp_icb_cmd_ready_511 = 1'b1;
  e603_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_delay_stage_511 (
    .i_vld(tmp_icb_cmd_valid_510), 
    .i_rdy(tmp_icb_cmd_ready_510), 
    .i_dat(tmp_icb_cmd_pack_510),
    .o_vld(tmp_icb_cmd_valid_511), 
    .o_rdy(delay_stage_select[511] ? byp_icb_cmd_ready : tmp_icb_cmd_ready_511), 
    .o_dat(tmp_icb_cmd_pack_511),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  assign byp_icb_cmd_valid      = 1'b0
                                | (tmp_icb_cmd_valid_0 & delay_stage_select[0])
                                | (tmp_icb_cmd_valid_1 & delay_stage_select[1])
                                | (tmp_icb_cmd_valid_2 & delay_stage_select[2])
                                | (tmp_icb_cmd_valid_3 & delay_stage_select[3])
                                | (tmp_icb_cmd_valid_4 & delay_stage_select[4])
                                | (tmp_icb_cmd_valid_5 & delay_stage_select[5])
                                | (tmp_icb_cmd_valid_6 & delay_stage_select[6])
                                | (tmp_icb_cmd_valid_7 & delay_stage_select[7])
                                | (tmp_icb_cmd_valid_8 & delay_stage_select[8])
                                | (tmp_icb_cmd_valid_9 & delay_stage_select[9])
                                | (tmp_icb_cmd_valid_10 & delay_stage_select[10])
                                | (tmp_icb_cmd_valid_11 & delay_stage_select[11])
                                | (tmp_icb_cmd_valid_12 & delay_stage_select[12])
                                | (tmp_icb_cmd_valid_13 & delay_stage_select[13])
                                | (tmp_icb_cmd_valid_14 & delay_stage_select[14])
                                | (tmp_icb_cmd_valid_15 & delay_stage_select[15])
                                | (tmp_icb_cmd_valid_16 & delay_stage_select[16])
                                | (tmp_icb_cmd_valid_17 & delay_stage_select[17])
                                | (tmp_icb_cmd_valid_18 & delay_stage_select[18])
                                | (tmp_icb_cmd_valid_19 & delay_stage_select[19])
                                | (tmp_icb_cmd_valid_20 & delay_stage_select[20])
                                | (tmp_icb_cmd_valid_21 & delay_stage_select[21])
                                | (tmp_icb_cmd_valid_22 & delay_stage_select[22])
                                | (tmp_icb_cmd_valid_23 & delay_stage_select[23])
                                | (tmp_icb_cmd_valid_24 & delay_stage_select[24])
                                | (tmp_icb_cmd_valid_25 & delay_stage_select[25])
                                | (tmp_icb_cmd_valid_26 & delay_stage_select[26])
                                | (tmp_icb_cmd_valid_27 & delay_stage_select[27])
                                | (tmp_icb_cmd_valid_28 & delay_stage_select[28])
                                | (tmp_icb_cmd_valid_29 & delay_stage_select[29])
                                | (tmp_icb_cmd_valid_30 & delay_stage_select[30])
                                | (tmp_icb_cmd_valid_31 & delay_stage_select[31])
                                | (tmp_icb_cmd_valid_32 & delay_stage_select[32])
                                | (tmp_icb_cmd_valid_33 & delay_stage_select[33])
                                | (tmp_icb_cmd_valid_34 & delay_stage_select[34])
                                | (tmp_icb_cmd_valid_35 & delay_stage_select[35])
                                | (tmp_icb_cmd_valid_36 & delay_stage_select[36])
                                | (tmp_icb_cmd_valid_37 & delay_stage_select[37])
                                | (tmp_icb_cmd_valid_38 & delay_stage_select[38])
                                | (tmp_icb_cmd_valid_39 & delay_stage_select[39])
                                | (tmp_icb_cmd_valid_40 & delay_stage_select[40])
                                | (tmp_icb_cmd_valid_41 & delay_stage_select[41])
                                | (tmp_icb_cmd_valid_42 & delay_stage_select[42])
                                | (tmp_icb_cmd_valid_43 & delay_stage_select[43])
                                | (tmp_icb_cmd_valid_44 & delay_stage_select[44])
                                | (tmp_icb_cmd_valid_45 & delay_stage_select[45])
                                | (tmp_icb_cmd_valid_46 & delay_stage_select[46])
                                | (tmp_icb_cmd_valid_47 & delay_stage_select[47])
                                | (tmp_icb_cmd_valid_48 & delay_stage_select[48])
                                | (tmp_icb_cmd_valid_49 & delay_stage_select[49])
                                | (tmp_icb_cmd_valid_50 & delay_stage_select[50])
                                | (tmp_icb_cmd_valid_51 & delay_stage_select[51])
                                | (tmp_icb_cmd_valid_52 & delay_stage_select[52])
                                | (tmp_icb_cmd_valid_53 & delay_stage_select[53])
                                | (tmp_icb_cmd_valid_54 & delay_stage_select[54])
                                | (tmp_icb_cmd_valid_55 & delay_stage_select[55])
                                | (tmp_icb_cmd_valid_56 & delay_stage_select[56])
                                | (tmp_icb_cmd_valid_57 & delay_stage_select[57])
                                | (tmp_icb_cmd_valid_58 & delay_stage_select[58])
                                | (tmp_icb_cmd_valid_59 & delay_stage_select[59])
                                | (tmp_icb_cmd_valid_60 & delay_stage_select[60])
                                | (tmp_icb_cmd_valid_61 & delay_stage_select[61])
                                | (tmp_icb_cmd_valid_62 & delay_stage_select[62])
                                | (tmp_icb_cmd_valid_63 & delay_stage_select[63])
                                | (tmp_icb_cmd_valid_64 & delay_stage_select[64])
                                | (tmp_icb_cmd_valid_65 & delay_stage_select[65])
                                | (tmp_icb_cmd_valid_66 & delay_stage_select[66])
                                | (tmp_icb_cmd_valid_67 & delay_stage_select[67])
                                | (tmp_icb_cmd_valid_68 & delay_stage_select[68])
                                | (tmp_icb_cmd_valid_69 & delay_stage_select[69])
                                | (tmp_icb_cmd_valid_70 & delay_stage_select[70])
                                | (tmp_icb_cmd_valid_71 & delay_stage_select[71])
                                | (tmp_icb_cmd_valid_72 & delay_stage_select[72])
                                | (tmp_icb_cmd_valid_73 & delay_stage_select[73])
                                | (tmp_icb_cmd_valid_74 & delay_stage_select[74])
                                | (tmp_icb_cmd_valid_75 & delay_stage_select[75])
                                | (tmp_icb_cmd_valid_76 & delay_stage_select[76])
                                | (tmp_icb_cmd_valid_77 & delay_stage_select[77])
                                | (tmp_icb_cmd_valid_78 & delay_stage_select[78])
                                | (tmp_icb_cmd_valid_79 & delay_stage_select[79])
                                | (tmp_icb_cmd_valid_80 & delay_stage_select[80])
                                | (tmp_icb_cmd_valid_81 & delay_stage_select[81])
                                | (tmp_icb_cmd_valid_82 & delay_stage_select[82])
                                | (tmp_icb_cmd_valid_83 & delay_stage_select[83])
                                | (tmp_icb_cmd_valid_84 & delay_stage_select[84])
                                | (tmp_icb_cmd_valid_85 & delay_stage_select[85])
                                | (tmp_icb_cmd_valid_86 & delay_stage_select[86])
                                | (tmp_icb_cmd_valid_87 & delay_stage_select[87])
                                | (tmp_icb_cmd_valid_88 & delay_stage_select[88])
                                | (tmp_icb_cmd_valid_89 & delay_stage_select[89])
                                | (tmp_icb_cmd_valid_90 & delay_stage_select[90])
                                | (tmp_icb_cmd_valid_91 & delay_stage_select[91])
                                | (tmp_icb_cmd_valid_92 & delay_stage_select[92])
                                | (tmp_icb_cmd_valid_93 & delay_stage_select[93])
                                | (tmp_icb_cmd_valid_94 & delay_stage_select[94])
                                | (tmp_icb_cmd_valid_95 & delay_stage_select[95])
                                | (tmp_icb_cmd_valid_96 & delay_stage_select[96])
                                | (tmp_icb_cmd_valid_97 & delay_stage_select[97])
                                | (tmp_icb_cmd_valid_98 & delay_stage_select[98])
                                | (tmp_icb_cmd_valid_99 & delay_stage_select[99])
                                | (tmp_icb_cmd_valid_100 & delay_stage_select[100])
                                | (tmp_icb_cmd_valid_101 & delay_stage_select[101])
                                | (tmp_icb_cmd_valid_102 & delay_stage_select[102])
                                | (tmp_icb_cmd_valid_103 & delay_stage_select[103])
                                | (tmp_icb_cmd_valid_104 & delay_stage_select[104])
                                | (tmp_icb_cmd_valid_105 & delay_stage_select[105])
                                | (tmp_icb_cmd_valid_106 & delay_stage_select[106])
                                | (tmp_icb_cmd_valid_107 & delay_stage_select[107])
                                | (tmp_icb_cmd_valid_108 & delay_stage_select[108])
                                | (tmp_icb_cmd_valid_109 & delay_stage_select[109])
                                | (tmp_icb_cmd_valid_110 & delay_stage_select[110])
                                | (tmp_icb_cmd_valid_111 & delay_stage_select[111])
                                | (tmp_icb_cmd_valid_112 & delay_stage_select[112])
                                | (tmp_icb_cmd_valid_113 & delay_stage_select[113])
                                | (tmp_icb_cmd_valid_114 & delay_stage_select[114])
                                | (tmp_icb_cmd_valid_115 & delay_stage_select[115])
                                | (tmp_icb_cmd_valid_116 & delay_stage_select[116])
                                | (tmp_icb_cmd_valid_117 & delay_stage_select[117])
                                | (tmp_icb_cmd_valid_118 & delay_stage_select[118])
                                | (tmp_icb_cmd_valid_119 & delay_stage_select[119])
                                | (tmp_icb_cmd_valid_120 & delay_stage_select[120])
                                | (tmp_icb_cmd_valid_121 & delay_stage_select[121])
                                | (tmp_icb_cmd_valid_122 & delay_stage_select[122])
                                | (tmp_icb_cmd_valid_123 & delay_stage_select[123])
                                | (tmp_icb_cmd_valid_124 & delay_stage_select[124])
                                | (tmp_icb_cmd_valid_125 & delay_stage_select[125])
                                | (tmp_icb_cmd_valid_126 & delay_stage_select[126])
                                | (tmp_icb_cmd_valid_127 & delay_stage_select[127])
                                | (tmp_icb_cmd_valid_128 & delay_stage_select[128])
                                | (tmp_icb_cmd_valid_129 & delay_stage_select[129])
                                | (tmp_icb_cmd_valid_130 & delay_stage_select[130])
                                | (tmp_icb_cmd_valid_131 & delay_stage_select[131])
                                | (tmp_icb_cmd_valid_132 & delay_stage_select[132])
                                | (tmp_icb_cmd_valid_133 & delay_stage_select[133])
                                | (tmp_icb_cmd_valid_134 & delay_stage_select[134])
                                | (tmp_icb_cmd_valid_135 & delay_stage_select[135])
                                | (tmp_icb_cmd_valid_136 & delay_stage_select[136])
                                | (tmp_icb_cmd_valid_137 & delay_stage_select[137])
                                | (tmp_icb_cmd_valid_138 & delay_stage_select[138])
                                | (tmp_icb_cmd_valid_139 & delay_stage_select[139])
                                | (tmp_icb_cmd_valid_140 & delay_stage_select[140])
                                | (tmp_icb_cmd_valid_141 & delay_stage_select[141])
                                | (tmp_icb_cmd_valid_142 & delay_stage_select[142])
                                | (tmp_icb_cmd_valid_143 & delay_stage_select[143])
                                | (tmp_icb_cmd_valid_144 & delay_stage_select[144])
                                | (tmp_icb_cmd_valid_145 & delay_stage_select[145])
                                | (tmp_icb_cmd_valid_146 & delay_stage_select[146])
                                | (tmp_icb_cmd_valid_147 & delay_stage_select[147])
                                | (tmp_icb_cmd_valid_148 & delay_stage_select[148])
                                | (tmp_icb_cmd_valid_149 & delay_stage_select[149])
                                | (tmp_icb_cmd_valid_150 & delay_stage_select[150])
                                | (tmp_icb_cmd_valid_151 & delay_stage_select[151])
                                | (tmp_icb_cmd_valid_152 & delay_stage_select[152])
                                | (tmp_icb_cmd_valid_153 & delay_stage_select[153])
                                | (tmp_icb_cmd_valid_154 & delay_stage_select[154])
                                | (tmp_icb_cmd_valid_155 & delay_stage_select[155])
                                | (tmp_icb_cmd_valid_156 & delay_stage_select[156])
                                | (tmp_icb_cmd_valid_157 & delay_stage_select[157])
                                | (tmp_icb_cmd_valid_158 & delay_stage_select[158])
                                | (tmp_icb_cmd_valid_159 & delay_stage_select[159])
                                | (tmp_icb_cmd_valid_160 & delay_stage_select[160])
                                | (tmp_icb_cmd_valid_161 & delay_stage_select[161])
                                | (tmp_icb_cmd_valid_162 & delay_stage_select[162])
                                | (tmp_icb_cmd_valid_163 & delay_stage_select[163])
                                | (tmp_icb_cmd_valid_164 & delay_stage_select[164])
                                | (tmp_icb_cmd_valid_165 & delay_stage_select[165])
                                | (tmp_icb_cmd_valid_166 & delay_stage_select[166])
                                | (tmp_icb_cmd_valid_167 & delay_stage_select[167])
                                | (tmp_icb_cmd_valid_168 & delay_stage_select[168])
                                | (tmp_icb_cmd_valid_169 & delay_stage_select[169])
                                | (tmp_icb_cmd_valid_170 & delay_stage_select[170])
                                | (tmp_icb_cmd_valid_171 & delay_stage_select[171])
                                | (tmp_icb_cmd_valid_172 & delay_stage_select[172])
                                | (tmp_icb_cmd_valid_173 & delay_stage_select[173])
                                | (tmp_icb_cmd_valid_174 & delay_stage_select[174])
                                | (tmp_icb_cmd_valid_175 & delay_stage_select[175])
                                | (tmp_icb_cmd_valid_176 & delay_stage_select[176])
                                | (tmp_icb_cmd_valid_177 & delay_stage_select[177])
                                | (tmp_icb_cmd_valid_178 & delay_stage_select[178])
                                | (tmp_icb_cmd_valid_179 & delay_stage_select[179])
                                | (tmp_icb_cmd_valid_180 & delay_stage_select[180])
                                | (tmp_icb_cmd_valid_181 & delay_stage_select[181])
                                | (tmp_icb_cmd_valid_182 & delay_stage_select[182])
                                | (tmp_icb_cmd_valid_183 & delay_stage_select[183])
                                | (tmp_icb_cmd_valid_184 & delay_stage_select[184])
                                | (tmp_icb_cmd_valid_185 & delay_stage_select[185])
                                | (tmp_icb_cmd_valid_186 & delay_stage_select[186])
                                | (tmp_icb_cmd_valid_187 & delay_stage_select[187])
                                | (tmp_icb_cmd_valid_188 & delay_stage_select[188])
                                | (tmp_icb_cmd_valid_189 & delay_stage_select[189])
                                | (tmp_icb_cmd_valid_190 & delay_stage_select[190])
                                | (tmp_icb_cmd_valid_191 & delay_stage_select[191])
                                | (tmp_icb_cmd_valid_192 & delay_stage_select[192])
                                | (tmp_icb_cmd_valid_193 & delay_stage_select[193])
                                | (tmp_icb_cmd_valid_194 & delay_stage_select[194])
                                | (tmp_icb_cmd_valid_195 & delay_stage_select[195])
                                | (tmp_icb_cmd_valid_196 & delay_stage_select[196])
                                | (tmp_icb_cmd_valid_197 & delay_stage_select[197])
                                | (tmp_icb_cmd_valid_198 & delay_stage_select[198])
                                | (tmp_icb_cmd_valid_199 & delay_stage_select[199])
                                | (tmp_icb_cmd_valid_200 & delay_stage_select[200])
                                | (tmp_icb_cmd_valid_201 & delay_stage_select[201])
                                | (tmp_icb_cmd_valid_202 & delay_stage_select[202])
                                | (tmp_icb_cmd_valid_203 & delay_stage_select[203])
                                | (tmp_icb_cmd_valid_204 & delay_stage_select[204])
                                | (tmp_icb_cmd_valid_205 & delay_stage_select[205])
                                | (tmp_icb_cmd_valid_206 & delay_stage_select[206])
                                | (tmp_icb_cmd_valid_207 & delay_stage_select[207])
                                | (tmp_icb_cmd_valid_208 & delay_stage_select[208])
                                | (tmp_icb_cmd_valid_209 & delay_stage_select[209])
                                | (tmp_icb_cmd_valid_210 & delay_stage_select[210])
                                | (tmp_icb_cmd_valid_211 & delay_stage_select[211])
                                | (tmp_icb_cmd_valid_212 & delay_stage_select[212])
                                | (tmp_icb_cmd_valid_213 & delay_stage_select[213])
                                | (tmp_icb_cmd_valid_214 & delay_stage_select[214])
                                | (tmp_icb_cmd_valid_215 & delay_stage_select[215])
                                | (tmp_icb_cmd_valid_216 & delay_stage_select[216])
                                | (tmp_icb_cmd_valid_217 & delay_stage_select[217])
                                | (tmp_icb_cmd_valid_218 & delay_stage_select[218])
                                | (tmp_icb_cmd_valid_219 & delay_stage_select[219])
                                | (tmp_icb_cmd_valid_220 & delay_stage_select[220])
                                | (tmp_icb_cmd_valid_221 & delay_stage_select[221])
                                | (tmp_icb_cmd_valid_222 & delay_stage_select[222])
                                | (tmp_icb_cmd_valid_223 & delay_stage_select[223])
                                | (tmp_icb_cmd_valid_224 & delay_stage_select[224])
                                | (tmp_icb_cmd_valid_225 & delay_stage_select[225])
                                | (tmp_icb_cmd_valid_226 & delay_stage_select[226])
                                | (tmp_icb_cmd_valid_227 & delay_stage_select[227])
                                | (tmp_icb_cmd_valid_228 & delay_stage_select[228])
                                | (tmp_icb_cmd_valid_229 & delay_stage_select[229])
                                | (tmp_icb_cmd_valid_230 & delay_stage_select[230])
                                | (tmp_icb_cmd_valid_231 & delay_stage_select[231])
                                | (tmp_icb_cmd_valid_232 & delay_stage_select[232])
                                | (tmp_icb_cmd_valid_233 & delay_stage_select[233])
                                | (tmp_icb_cmd_valid_234 & delay_stage_select[234])
                                | (tmp_icb_cmd_valid_235 & delay_stage_select[235])
                                | (tmp_icb_cmd_valid_236 & delay_stage_select[236])
                                | (tmp_icb_cmd_valid_237 & delay_stage_select[237])
                                | (tmp_icb_cmd_valid_238 & delay_stage_select[238])
                                | (tmp_icb_cmd_valid_239 & delay_stage_select[239])
                                | (tmp_icb_cmd_valid_240 & delay_stage_select[240])
                                | (tmp_icb_cmd_valid_241 & delay_stage_select[241])
                                | (tmp_icb_cmd_valid_242 & delay_stage_select[242])
                                | (tmp_icb_cmd_valid_243 & delay_stage_select[243])
                                | (tmp_icb_cmd_valid_244 & delay_stage_select[244])
                                | (tmp_icb_cmd_valid_245 & delay_stage_select[245])
                                | (tmp_icb_cmd_valid_246 & delay_stage_select[246])
                                | (tmp_icb_cmd_valid_247 & delay_stage_select[247])
                                | (tmp_icb_cmd_valid_248 & delay_stage_select[248])
                                | (tmp_icb_cmd_valid_249 & delay_stage_select[249])
                                | (tmp_icb_cmd_valid_250 & delay_stage_select[250])
                                | (tmp_icb_cmd_valid_251 & delay_stage_select[251])
                                | (tmp_icb_cmd_valid_252 & delay_stage_select[252])
                                | (tmp_icb_cmd_valid_253 & delay_stage_select[253])
                                | (tmp_icb_cmd_valid_254 & delay_stage_select[254])
                                | (tmp_icb_cmd_valid_255 & delay_stage_select[255])
                                | (tmp_icb_cmd_valid_256 & delay_stage_select[256])
                                | (tmp_icb_cmd_valid_257 & delay_stage_select[257])
                                | (tmp_icb_cmd_valid_258 & delay_stage_select[258])
                                | (tmp_icb_cmd_valid_259 & delay_stage_select[259])
                                | (tmp_icb_cmd_valid_260 & delay_stage_select[260])
                                | (tmp_icb_cmd_valid_261 & delay_stage_select[261])
                                | (tmp_icb_cmd_valid_262 & delay_stage_select[262])
                                | (tmp_icb_cmd_valid_263 & delay_stage_select[263])
                                | (tmp_icb_cmd_valid_264 & delay_stage_select[264])
                                | (tmp_icb_cmd_valid_265 & delay_stage_select[265])
                                | (tmp_icb_cmd_valid_266 & delay_stage_select[266])
                                | (tmp_icb_cmd_valid_267 & delay_stage_select[267])
                                | (tmp_icb_cmd_valid_268 & delay_stage_select[268])
                                | (tmp_icb_cmd_valid_269 & delay_stage_select[269])
                                | (tmp_icb_cmd_valid_270 & delay_stage_select[270])
                                | (tmp_icb_cmd_valid_271 & delay_stage_select[271])
                                | (tmp_icb_cmd_valid_272 & delay_stage_select[272])
                                | (tmp_icb_cmd_valid_273 & delay_stage_select[273])
                                | (tmp_icb_cmd_valid_274 & delay_stage_select[274])
                                | (tmp_icb_cmd_valid_275 & delay_stage_select[275])
                                | (tmp_icb_cmd_valid_276 & delay_stage_select[276])
                                | (tmp_icb_cmd_valid_277 & delay_stage_select[277])
                                | (tmp_icb_cmd_valid_278 & delay_stage_select[278])
                                | (tmp_icb_cmd_valid_279 & delay_stage_select[279])
                                | (tmp_icb_cmd_valid_280 & delay_stage_select[280])
                                | (tmp_icb_cmd_valid_281 & delay_stage_select[281])
                                | (tmp_icb_cmd_valid_282 & delay_stage_select[282])
                                | (tmp_icb_cmd_valid_283 & delay_stage_select[283])
                                | (tmp_icb_cmd_valid_284 & delay_stage_select[284])
                                | (tmp_icb_cmd_valid_285 & delay_stage_select[285])
                                | (tmp_icb_cmd_valid_286 & delay_stage_select[286])
                                | (tmp_icb_cmd_valid_287 & delay_stage_select[287])
                                | (tmp_icb_cmd_valid_288 & delay_stage_select[288])
                                | (tmp_icb_cmd_valid_289 & delay_stage_select[289])
                                | (tmp_icb_cmd_valid_290 & delay_stage_select[290])
                                | (tmp_icb_cmd_valid_291 & delay_stage_select[291])
                                | (tmp_icb_cmd_valid_292 & delay_stage_select[292])
                                | (tmp_icb_cmd_valid_293 & delay_stage_select[293])
                                | (tmp_icb_cmd_valid_294 & delay_stage_select[294])
                                | (tmp_icb_cmd_valid_295 & delay_stage_select[295])
                                | (tmp_icb_cmd_valid_296 & delay_stage_select[296])
                                | (tmp_icb_cmd_valid_297 & delay_stage_select[297])
                                | (tmp_icb_cmd_valid_298 & delay_stage_select[298])
                                | (tmp_icb_cmd_valid_299 & delay_stage_select[299])
                                | (tmp_icb_cmd_valid_300 & delay_stage_select[300])
                                | (tmp_icb_cmd_valid_301 & delay_stage_select[301])
                                | (tmp_icb_cmd_valid_302 & delay_stage_select[302])
                                | (tmp_icb_cmd_valid_303 & delay_stage_select[303])
                                | (tmp_icb_cmd_valid_304 & delay_stage_select[304])
                                | (tmp_icb_cmd_valid_305 & delay_stage_select[305])
                                | (tmp_icb_cmd_valid_306 & delay_stage_select[306])
                                | (tmp_icb_cmd_valid_307 & delay_stage_select[307])
                                | (tmp_icb_cmd_valid_308 & delay_stage_select[308])
                                | (tmp_icb_cmd_valid_309 & delay_stage_select[309])
                                | (tmp_icb_cmd_valid_310 & delay_stage_select[310])
                                | (tmp_icb_cmd_valid_311 & delay_stage_select[311])
                                | (tmp_icb_cmd_valid_312 & delay_stage_select[312])
                                | (tmp_icb_cmd_valid_313 & delay_stage_select[313])
                                | (tmp_icb_cmd_valid_314 & delay_stage_select[314])
                                | (tmp_icb_cmd_valid_315 & delay_stage_select[315])
                                | (tmp_icb_cmd_valid_316 & delay_stage_select[316])
                                | (tmp_icb_cmd_valid_317 & delay_stage_select[317])
                                | (tmp_icb_cmd_valid_318 & delay_stage_select[318])
                                | (tmp_icb_cmd_valid_319 & delay_stage_select[319])
                                | (tmp_icb_cmd_valid_320 & delay_stage_select[320])
                                | (tmp_icb_cmd_valid_321 & delay_stage_select[321])
                                | (tmp_icb_cmd_valid_322 & delay_stage_select[322])
                                | (tmp_icb_cmd_valid_323 & delay_stage_select[323])
                                | (tmp_icb_cmd_valid_324 & delay_stage_select[324])
                                | (tmp_icb_cmd_valid_325 & delay_stage_select[325])
                                | (tmp_icb_cmd_valid_326 & delay_stage_select[326])
                                | (tmp_icb_cmd_valid_327 & delay_stage_select[327])
                                | (tmp_icb_cmd_valid_328 & delay_stage_select[328])
                                | (tmp_icb_cmd_valid_329 & delay_stage_select[329])
                                | (tmp_icb_cmd_valid_330 & delay_stage_select[330])
                                | (tmp_icb_cmd_valid_331 & delay_stage_select[331])
                                | (tmp_icb_cmd_valid_332 & delay_stage_select[332])
                                | (tmp_icb_cmd_valid_333 & delay_stage_select[333])
                                | (tmp_icb_cmd_valid_334 & delay_stage_select[334])
                                | (tmp_icb_cmd_valid_335 & delay_stage_select[335])
                                | (tmp_icb_cmd_valid_336 & delay_stage_select[336])
                                | (tmp_icb_cmd_valid_337 & delay_stage_select[337])
                                | (tmp_icb_cmd_valid_338 & delay_stage_select[338])
                                | (tmp_icb_cmd_valid_339 & delay_stage_select[339])
                                | (tmp_icb_cmd_valid_340 & delay_stage_select[340])
                                | (tmp_icb_cmd_valid_341 & delay_stage_select[341])
                                | (tmp_icb_cmd_valid_342 & delay_stage_select[342])
                                | (tmp_icb_cmd_valid_343 & delay_stage_select[343])
                                | (tmp_icb_cmd_valid_344 & delay_stage_select[344])
                                | (tmp_icb_cmd_valid_345 & delay_stage_select[345])
                                | (tmp_icb_cmd_valid_346 & delay_stage_select[346])
                                | (tmp_icb_cmd_valid_347 & delay_stage_select[347])
                                | (tmp_icb_cmd_valid_348 & delay_stage_select[348])
                                | (tmp_icb_cmd_valid_349 & delay_stage_select[349])
                                | (tmp_icb_cmd_valid_350 & delay_stage_select[350])
                                | (tmp_icb_cmd_valid_351 & delay_stage_select[351])
                                | (tmp_icb_cmd_valid_352 & delay_stage_select[352])
                                | (tmp_icb_cmd_valid_353 & delay_stage_select[353])
                                | (tmp_icb_cmd_valid_354 & delay_stage_select[354])
                                | (tmp_icb_cmd_valid_355 & delay_stage_select[355])
                                | (tmp_icb_cmd_valid_356 & delay_stage_select[356])
                                | (tmp_icb_cmd_valid_357 & delay_stage_select[357])
                                | (tmp_icb_cmd_valid_358 & delay_stage_select[358])
                                | (tmp_icb_cmd_valid_359 & delay_stage_select[359])
                                | (tmp_icb_cmd_valid_360 & delay_stage_select[360])
                                | (tmp_icb_cmd_valid_361 & delay_stage_select[361])
                                | (tmp_icb_cmd_valid_362 & delay_stage_select[362])
                                | (tmp_icb_cmd_valid_363 & delay_stage_select[363])
                                | (tmp_icb_cmd_valid_364 & delay_stage_select[364])
                                | (tmp_icb_cmd_valid_365 & delay_stage_select[365])
                                | (tmp_icb_cmd_valid_366 & delay_stage_select[366])
                                | (tmp_icb_cmd_valid_367 & delay_stage_select[367])
                                | (tmp_icb_cmd_valid_368 & delay_stage_select[368])
                                | (tmp_icb_cmd_valid_369 & delay_stage_select[369])
                                | (tmp_icb_cmd_valid_370 & delay_stage_select[370])
                                | (tmp_icb_cmd_valid_371 & delay_stage_select[371])
                                | (tmp_icb_cmd_valid_372 & delay_stage_select[372])
                                | (tmp_icb_cmd_valid_373 & delay_stage_select[373])
                                | (tmp_icb_cmd_valid_374 & delay_stage_select[374])
                                | (tmp_icb_cmd_valid_375 & delay_stage_select[375])
                                | (tmp_icb_cmd_valid_376 & delay_stage_select[376])
                                | (tmp_icb_cmd_valid_377 & delay_stage_select[377])
                                | (tmp_icb_cmd_valid_378 & delay_stage_select[378])
                                | (tmp_icb_cmd_valid_379 & delay_stage_select[379])
                                | (tmp_icb_cmd_valid_380 & delay_stage_select[380])
                                | (tmp_icb_cmd_valid_381 & delay_stage_select[381])
                                | (tmp_icb_cmd_valid_382 & delay_stage_select[382])
                                | (tmp_icb_cmd_valid_383 & delay_stage_select[383])
                                | (tmp_icb_cmd_valid_384 & delay_stage_select[384])
                                | (tmp_icb_cmd_valid_385 & delay_stage_select[385])
                                | (tmp_icb_cmd_valid_386 & delay_stage_select[386])
                                | (tmp_icb_cmd_valid_387 & delay_stage_select[387])
                                | (tmp_icb_cmd_valid_388 & delay_stage_select[388])
                                | (tmp_icb_cmd_valid_389 & delay_stage_select[389])
                                | (tmp_icb_cmd_valid_390 & delay_stage_select[390])
                                | (tmp_icb_cmd_valid_391 & delay_stage_select[391])
                                | (tmp_icb_cmd_valid_392 & delay_stage_select[392])
                                | (tmp_icb_cmd_valid_393 & delay_stage_select[393])
                                | (tmp_icb_cmd_valid_394 & delay_stage_select[394])
                                | (tmp_icb_cmd_valid_395 & delay_stage_select[395])
                                | (tmp_icb_cmd_valid_396 & delay_stage_select[396])
                                | (tmp_icb_cmd_valid_397 & delay_stage_select[397])
                                | (tmp_icb_cmd_valid_398 & delay_stage_select[398])
                                | (tmp_icb_cmd_valid_399 & delay_stage_select[399])
                                | (tmp_icb_cmd_valid_400 & delay_stage_select[400])
                                | (tmp_icb_cmd_valid_401 & delay_stage_select[401])
                                | (tmp_icb_cmd_valid_402 & delay_stage_select[402])
                                | (tmp_icb_cmd_valid_403 & delay_stage_select[403])
                                | (tmp_icb_cmd_valid_404 & delay_stage_select[404])
                                | (tmp_icb_cmd_valid_405 & delay_stage_select[405])
                                | (tmp_icb_cmd_valid_406 & delay_stage_select[406])
                                | (tmp_icb_cmd_valid_407 & delay_stage_select[407])
                                | (tmp_icb_cmd_valid_408 & delay_stage_select[408])
                                | (tmp_icb_cmd_valid_409 & delay_stage_select[409])
                                | (tmp_icb_cmd_valid_410 & delay_stage_select[410])
                                | (tmp_icb_cmd_valid_411 & delay_stage_select[411])
                                | (tmp_icb_cmd_valid_412 & delay_stage_select[412])
                                | (tmp_icb_cmd_valid_413 & delay_stage_select[413])
                                | (tmp_icb_cmd_valid_414 & delay_stage_select[414])
                                | (tmp_icb_cmd_valid_415 & delay_stage_select[415])
                                | (tmp_icb_cmd_valid_416 & delay_stage_select[416])
                                | (tmp_icb_cmd_valid_417 & delay_stage_select[417])
                                | (tmp_icb_cmd_valid_418 & delay_stage_select[418])
                                | (tmp_icb_cmd_valid_419 & delay_stage_select[419])
                                | (tmp_icb_cmd_valid_420 & delay_stage_select[420])
                                | (tmp_icb_cmd_valid_421 & delay_stage_select[421])
                                | (tmp_icb_cmd_valid_422 & delay_stage_select[422])
                                | (tmp_icb_cmd_valid_423 & delay_stage_select[423])
                                | (tmp_icb_cmd_valid_424 & delay_stage_select[424])
                                | (tmp_icb_cmd_valid_425 & delay_stage_select[425])
                                | (tmp_icb_cmd_valid_426 & delay_stage_select[426])
                                | (tmp_icb_cmd_valid_427 & delay_stage_select[427])
                                | (tmp_icb_cmd_valid_428 & delay_stage_select[428])
                                | (tmp_icb_cmd_valid_429 & delay_stage_select[429])
                                | (tmp_icb_cmd_valid_430 & delay_stage_select[430])
                                | (tmp_icb_cmd_valid_431 & delay_stage_select[431])
                                | (tmp_icb_cmd_valid_432 & delay_stage_select[432])
                                | (tmp_icb_cmd_valid_433 & delay_stage_select[433])
                                | (tmp_icb_cmd_valid_434 & delay_stage_select[434])
                                | (tmp_icb_cmd_valid_435 & delay_stage_select[435])
                                | (tmp_icb_cmd_valid_436 & delay_stage_select[436])
                                | (tmp_icb_cmd_valid_437 & delay_stage_select[437])
                                | (tmp_icb_cmd_valid_438 & delay_stage_select[438])
                                | (tmp_icb_cmd_valid_439 & delay_stage_select[439])
                                | (tmp_icb_cmd_valid_440 & delay_stage_select[440])
                                | (tmp_icb_cmd_valid_441 & delay_stage_select[441])
                                | (tmp_icb_cmd_valid_442 & delay_stage_select[442])
                                | (tmp_icb_cmd_valid_443 & delay_stage_select[443])
                                | (tmp_icb_cmd_valid_444 & delay_stage_select[444])
                                | (tmp_icb_cmd_valid_445 & delay_stage_select[445])
                                | (tmp_icb_cmd_valid_446 & delay_stage_select[446])
                                | (tmp_icb_cmd_valid_447 & delay_stage_select[447])
                                | (tmp_icb_cmd_valid_448 & delay_stage_select[448])
                                | (tmp_icb_cmd_valid_449 & delay_stage_select[449])
                                | (tmp_icb_cmd_valid_450 & delay_stage_select[450])
                                | (tmp_icb_cmd_valid_451 & delay_stage_select[451])
                                | (tmp_icb_cmd_valid_452 & delay_stage_select[452])
                                | (tmp_icb_cmd_valid_453 & delay_stage_select[453])
                                | (tmp_icb_cmd_valid_454 & delay_stage_select[454])
                                | (tmp_icb_cmd_valid_455 & delay_stage_select[455])
                                | (tmp_icb_cmd_valid_456 & delay_stage_select[456])
                                | (tmp_icb_cmd_valid_457 & delay_stage_select[457])
                                | (tmp_icb_cmd_valid_458 & delay_stage_select[458])
                                | (tmp_icb_cmd_valid_459 & delay_stage_select[459])
                                | (tmp_icb_cmd_valid_460 & delay_stage_select[460])
                                | (tmp_icb_cmd_valid_461 & delay_stage_select[461])
                                | (tmp_icb_cmd_valid_462 & delay_stage_select[462])
                                | (tmp_icb_cmd_valid_463 & delay_stage_select[463])
                                | (tmp_icb_cmd_valid_464 & delay_stage_select[464])
                                | (tmp_icb_cmd_valid_465 & delay_stage_select[465])
                                | (tmp_icb_cmd_valid_466 & delay_stage_select[466])
                                | (tmp_icb_cmd_valid_467 & delay_stage_select[467])
                                | (tmp_icb_cmd_valid_468 & delay_stage_select[468])
                                | (tmp_icb_cmd_valid_469 & delay_stage_select[469])
                                | (tmp_icb_cmd_valid_470 & delay_stage_select[470])
                                | (tmp_icb_cmd_valid_471 & delay_stage_select[471])
                                | (tmp_icb_cmd_valid_472 & delay_stage_select[472])
                                | (tmp_icb_cmd_valid_473 & delay_stage_select[473])
                                | (tmp_icb_cmd_valid_474 & delay_stage_select[474])
                                | (tmp_icb_cmd_valid_475 & delay_stage_select[475])
                                | (tmp_icb_cmd_valid_476 & delay_stage_select[476])
                                | (tmp_icb_cmd_valid_477 & delay_stage_select[477])
                                | (tmp_icb_cmd_valid_478 & delay_stage_select[478])
                                | (tmp_icb_cmd_valid_479 & delay_stage_select[479])
                                | (tmp_icb_cmd_valid_480 & delay_stage_select[480])
                                | (tmp_icb_cmd_valid_481 & delay_stage_select[481])
                                | (tmp_icb_cmd_valid_482 & delay_stage_select[482])
                                | (tmp_icb_cmd_valid_483 & delay_stage_select[483])
                                | (tmp_icb_cmd_valid_484 & delay_stage_select[484])
                                | (tmp_icb_cmd_valid_485 & delay_stage_select[485])
                                | (tmp_icb_cmd_valid_486 & delay_stage_select[486])
                                | (tmp_icb_cmd_valid_487 & delay_stage_select[487])
                                | (tmp_icb_cmd_valid_488 & delay_stage_select[488])
                                | (tmp_icb_cmd_valid_489 & delay_stage_select[489])
                                | (tmp_icb_cmd_valid_490 & delay_stage_select[490])
                                | (tmp_icb_cmd_valid_491 & delay_stage_select[491])
                                | (tmp_icb_cmd_valid_492 & delay_stage_select[492])
                                | (tmp_icb_cmd_valid_493 & delay_stage_select[493])
                                | (tmp_icb_cmd_valid_494 & delay_stage_select[494])
                                | (tmp_icb_cmd_valid_495 & delay_stage_select[495])
                                | (tmp_icb_cmd_valid_496 & delay_stage_select[496])
                                | (tmp_icb_cmd_valid_497 & delay_stage_select[497])
                                | (tmp_icb_cmd_valid_498 & delay_stage_select[498])
                                | (tmp_icb_cmd_valid_499 & delay_stage_select[499])
                                | (tmp_icb_cmd_valid_500 & delay_stage_select[500])
                                | (tmp_icb_cmd_valid_501 & delay_stage_select[501])
                                | (tmp_icb_cmd_valid_502 & delay_stage_select[502])
                                | (tmp_icb_cmd_valid_503 & delay_stage_select[503])
                                | (tmp_icb_cmd_valid_504 & delay_stage_select[504])
                                | (tmp_icb_cmd_valid_505 & delay_stage_select[505])
                                | (tmp_icb_cmd_valid_506 & delay_stage_select[506])
                                | (tmp_icb_cmd_valid_507 & delay_stage_select[507])
                                | (tmp_icb_cmd_valid_508 & delay_stage_select[508])
                                | (tmp_icb_cmd_valid_509 & delay_stage_select[509])
                                | (tmp_icb_cmd_valid_510 & delay_stage_select[510])
                                | (tmp_icb_cmd_valid_511 & delay_stage_select[511])
                                ;
  assign byp_icb_cmd_o_pack     = {BUF_CMD_PACK_W{1'b0}}
                                | (tmp_icb_cmd_pack_0 & {BUF_CMD_PACK_W{delay_stage_select[0]}})
                                | (tmp_icb_cmd_pack_1 & {BUF_CMD_PACK_W{delay_stage_select[1]}})
                                | (tmp_icb_cmd_pack_2 & {BUF_CMD_PACK_W{delay_stage_select[2]}})
                                | (tmp_icb_cmd_pack_3 & {BUF_CMD_PACK_W{delay_stage_select[3]}})
                                | (tmp_icb_cmd_pack_4 & {BUF_CMD_PACK_W{delay_stage_select[4]}})
                                | (tmp_icb_cmd_pack_5 & {BUF_CMD_PACK_W{delay_stage_select[5]}})
                                | (tmp_icb_cmd_pack_6 & {BUF_CMD_PACK_W{delay_stage_select[6]}})
                                | (tmp_icb_cmd_pack_7 & {BUF_CMD_PACK_W{delay_stage_select[7]}})
                                | (tmp_icb_cmd_pack_8 & {BUF_CMD_PACK_W{delay_stage_select[8]}})
                                | (tmp_icb_cmd_pack_9 & {BUF_CMD_PACK_W{delay_stage_select[9]}})
                                | (tmp_icb_cmd_pack_10 & {BUF_CMD_PACK_W{delay_stage_select[10]}})
                                | (tmp_icb_cmd_pack_11 & {BUF_CMD_PACK_W{delay_stage_select[11]}})
                                | (tmp_icb_cmd_pack_12 & {BUF_CMD_PACK_W{delay_stage_select[12]}})
                                | (tmp_icb_cmd_pack_13 & {BUF_CMD_PACK_W{delay_stage_select[13]}})
                                | (tmp_icb_cmd_pack_14 & {BUF_CMD_PACK_W{delay_stage_select[14]}})
                                | (tmp_icb_cmd_pack_15 & {BUF_CMD_PACK_W{delay_stage_select[15]}})
                                | (tmp_icb_cmd_pack_16 & {BUF_CMD_PACK_W{delay_stage_select[16]}})
                                | (tmp_icb_cmd_pack_17 & {BUF_CMD_PACK_W{delay_stage_select[17]}})
                                | (tmp_icb_cmd_pack_18 & {BUF_CMD_PACK_W{delay_stage_select[18]}})
                                | (tmp_icb_cmd_pack_19 & {BUF_CMD_PACK_W{delay_stage_select[19]}})
                                | (tmp_icb_cmd_pack_20 & {BUF_CMD_PACK_W{delay_stage_select[20]}})
                                | (tmp_icb_cmd_pack_21 & {BUF_CMD_PACK_W{delay_stage_select[21]}})
                                | (tmp_icb_cmd_pack_22 & {BUF_CMD_PACK_W{delay_stage_select[22]}})
                                | (tmp_icb_cmd_pack_23 & {BUF_CMD_PACK_W{delay_stage_select[23]}})
                                | (tmp_icb_cmd_pack_24 & {BUF_CMD_PACK_W{delay_stage_select[24]}})
                                | (tmp_icb_cmd_pack_25 & {BUF_CMD_PACK_W{delay_stage_select[25]}})
                                | (tmp_icb_cmd_pack_26 & {BUF_CMD_PACK_W{delay_stage_select[26]}})
                                | (tmp_icb_cmd_pack_27 & {BUF_CMD_PACK_W{delay_stage_select[27]}})
                                | (tmp_icb_cmd_pack_28 & {BUF_CMD_PACK_W{delay_stage_select[28]}})
                                | (tmp_icb_cmd_pack_29 & {BUF_CMD_PACK_W{delay_stage_select[29]}})
                                | (tmp_icb_cmd_pack_30 & {BUF_CMD_PACK_W{delay_stage_select[30]}})
                                | (tmp_icb_cmd_pack_31 & {BUF_CMD_PACK_W{delay_stage_select[31]}})
                                | (tmp_icb_cmd_pack_32 & {BUF_CMD_PACK_W{delay_stage_select[32]}})
                                | (tmp_icb_cmd_pack_33 & {BUF_CMD_PACK_W{delay_stage_select[33]}})
                                | (tmp_icb_cmd_pack_34 & {BUF_CMD_PACK_W{delay_stage_select[34]}})
                                | (tmp_icb_cmd_pack_35 & {BUF_CMD_PACK_W{delay_stage_select[35]}})
                                | (tmp_icb_cmd_pack_36 & {BUF_CMD_PACK_W{delay_stage_select[36]}})
                                | (tmp_icb_cmd_pack_37 & {BUF_CMD_PACK_W{delay_stage_select[37]}})
                                | (tmp_icb_cmd_pack_38 & {BUF_CMD_PACK_W{delay_stage_select[38]}})
                                | (tmp_icb_cmd_pack_39 & {BUF_CMD_PACK_W{delay_stage_select[39]}})
                                | (tmp_icb_cmd_pack_40 & {BUF_CMD_PACK_W{delay_stage_select[40]}})
                                | (tmp_icb_cmd_pack_41 & {BUF_CMD_PACK_W{delay_stage_select[41]}})
                                | (tmp_icb_cmd_pack_42 & {BUF_CMD_PACK_W{delay_stage_select[42]}})
                                | (tmp_icb_cmd_pack_43 & {BUF_CMD_PACK_W{delay_stage_select[43]}})
                                | (tmp_icb_cmd_pack_44 & {BUF_CMD_PACK_W{delay_stage_select[44]}})
                                | (tmp_icb_cmd_pack_45 & {BUF_CMD_PACK_W{delay_stage_select[45]}})
                                | (tmp_icb_cmd_pack_46 & {BUF_CMD_PACK_W{delay_stage_select[46]}})
                                | (tmp_icb_cmd_pack_47 & {BUF_CMD_PACK_W{delay_stage_select[47]}})
                                | (tmp_icb_cmd_pack_48 & {BUF_CMD_PACK_W{delay_stage_select[48]}})
                                | (tmp_icb_cmd_pack_49 & {BUF_CMD_PACK_W{delay_stage_select[49]}})
                                | (tmp_icb_cmd_pack_50 & {BUF_CMD_PACK_W{delay_stage_select[50]}})
                                | (tmp_icb_cmd_pack_51 & {BUF_CMD_PACK_W{delay_stage_select[51]}})
                                | (tmp_icb_cmd_pack_52 & {BUF_CMD_PACK_W{delay_stage_select[52]}})
                                | (tmp_icb_cmd_pack_53 & {BUF_CMD_PACK_W{delay_stage_select[53]}})
                                | (tmp_icb_cmd_pack_54 & {BUF_CMD_PACK_W{delay_stage_select[54]}})
                                | (tmp_icb_cmd_pack_55 & {BUF_CMD_PACK_W{delay_stage_select[55]}})
                                | (tmp_icb_cmd_pack_56 & {BUF_CMD_PACK_W{delay_stage_select[56]}})
                                | (tmp_icb_cmd_pack_57 & {BUF_CMD_PACK_W{delay_stage_select[57]}})
                                | (tmp_icb_cmd_pack_58 & {BUF_CMD_PACK_W{delay_stage_select[58]}})
                                | (tmp_icb_cmd_pack_59 & {BUF_CMD_PACK_W{delay_stage_select[59]}})
                                | (tmp_icb_cmd_pack_60 & {BUF_CMD_PACK_W{delay_stage_select[60]}})
                                | (tmp_icb_cmd_pack_61 & {BUF_CMD_PACK_W{delay_stage_select[61]}})
                                | (tmp_icb_cmd_pack_62 & {BUF_CMD_PACK_W{delay_stage_select[62]}})
                                | (tmp_icb_cmd_pack_63 & {BUF_CMD_PACK_W{delay_stage_select[63]}})
                                | (tmp_icb_cmd_pack_64 & {BUF_CMD_PACK_W{delay_stage_select[64]}})
                                | (tmp_icb_cmd_pack_65 & {BUF_CMD_PACK_W{delay_stage_select[65]}})
                                | (tmp_icb_cmd_pack_66 & {BUF_CMD_PACK_W{delay_stage_select[66]}})
                                | (tmp_icb_cmd_pack_67 & {BUF_CMD_PACK_W{delay_stage_select[67]}})
                                | (tmp_icb_cmd_pack_68 & {BUF_CMD_PACK_W{delay_stage_select[68]}})
                                | (tmp_icb_cmd_pack_69 & {BUF_CMD_PACK_W{delay_stage_select[69]}})
                                | (tmp_icb_cmd_pack_70 & {BUF_CMD_PACK_W{delay_stage_select[70]}})
                                | (tmp_icb_cmd_pack_71 & {BUF_CMD_PACK_W{delay_stage_select[71]}})
                                | (tmp_icb_cmd_pack_72 & {BUF_CMD_PACK_W{delay_stage_select[72]}})
                                | (tmp_icb_cmd_pack_73 & {BUF_CMD_PACK_W{delay_stage_select[73]}})
                                | (tmp_icb_cmd_pack_74 & {BUF_CMD_PACK_W{delay_stage_select[74]}})
                                | (tmp_icb_cmd_pack_75 & {BUF_CMD_PACK_W{delay_stage_select[75]}})
                                | (tmp_icb_cmd_pack_76 & {BUF_CMD_PACK_W{delay_stage_select[76]}})
                                | (tmp_icb_cmd_pack_77 & {BUF_CMD_PACK_W{delay_stage_select[77]}})
                                | (tmp_icb_cmd_pack_78 & {BUF_CMD_PACK_W{delay_stage_select[78]}})
                                | (tmp_icb_cmd_pack_79 & {BUF_CMD_PACK_W{delay_stage_select[79]}})
                                | (tmp_icb_cmd_pack_80 & {BUF_CMD_PACK_W{delay_stage_select[80]}})
                                | (tmp_icb_cmd_pack_81 & {BUF_CMD_PACK_W{delay_stage_select[81]}})
                                | (tmp_icb_cmd_pack_82 & {BUF_CMD_PACK_W{delay_stage_select[82]}})
                                | (tmp_icb_cmd_pack_83 & {BUF_CMD_PACK_W{delay_stage_select[83]}})
                                | (tmp_icb_cmd_pack_84 & {BUF_CMD_PACK_W{delay_stage_select[84]}})
                                | (tmp_icb_cmd_pack_85 & {BUF_CMD_PACK_W{delay_stage_select[85]}})
                                | (tmp_icb_cmd_pack_86 & {BUF_CMD_PACK_W{delay_stage_select[86]}})
                                | (tmp_icb_cmd_pack_87 & {BUF_CMD_PACK_W{delay_stage_select[87]}})
                                | (tmp_icb_cmd_pack_88 & {BUF_CMD_PACK_W{delay_stage_select[88]}})
                                | (tmp_icb_cmd_pack_89 & {BUF_CMD_PACK_W{delay_stage_select[89]}})
                                | (tmp_icb_cmd_pack_90 & {BUF_CMD_PACK_W{delay_stage_select[90]}})
                                | (tmp_icb_cmd_pack_91 & {BUF_CMD_PACK_W{delay_stage_select[91]}})
                                | (tmp_icb_cmd_pack_92 & {BUF_CMD_PACK_W{delay_stage_select[92]}})
                                | (tmp_icb_cmd_pack_93 & {BUF_CMD_PACK_W{delay_stage_select[93]}})
                                | (tmp_icb_cmd_pack_94 & {BUF_CMD_PACK_W{delay_stage_select[94]}})
                                | (tmp_icb_cmd_pack_95 & {BUF_CMD_PACK_W{delay_stage_select[95]}})
                                | (tmp_icb_cmd_pack_96 & {BUF_CMD_PACK_W{delay_stage_select[96]}})
                                | (tmp_icb_cmd_pack_97 & {BUF_CMD_PACK_W{delay_stage_select[97]}})
                                | (tmp_icb_cmd_pack_98 & {BUF_CMD_PACK_W{delay_stage_select[98]}})
                                | (tmp_icb_cmd_pack_99 & {BUF_CMD_PACK_W{delay_stage_select[99]}})
                                | (tmp_icb_cmd_pack_100 & {BUF_CMD_PACK_W{delay_stage_select[100]}})
                                | (tmp_icb_cmd_pack_101 & {BUF_CMD_PACK_W{delay_stage_select[101]}})
                                | (tmp_icb_cmd_pack_102 & {BUF_CMD_PACK_W{delay_stage_select[102]}})
                                | (tmp_icb_cmd_pack_103 & {BUF_CMD_PACK_W{delay_stage_select[103]}})
                                | (tmp_icb_cmd_pack_104 & {BUF_CMD_PACK_W{delay_stage_select[104]}})
                                | (tmp_icb_cmd_pack_105 & {BUF_CMD_PACK_W{delay_stage_select[105]}})
                                | (tmp_icb_cmd_pack_106 & {BUF_CMD_PACK_W{delay_stage_select[106]}})
                                | (tmp_icb_cmd_pack_107 & {BUF_CMD_PACK_W{delay_stage_select[107]}})
                                | (tmp_icb_cmd_pack_108 & {BUF_CMD_PACK_W{delay_stage_select[108]}})
                                | (tmp_icb_cmd_pack_109 & {BUF_CMD_PACK_W{delay_stage_select[109]}})
                                | (tmp_icb_cmd_pack_110 & {BUF_CMD_PACK_W{delay_stage_select[110]}})
                                | (tmp_icb_cmd_pack_111 & {BUF_CMD_PACK_W{delay_stage_select[111]}})
                                | (tmp_icb_cmd_pack_112 & {BUF_CMD_PACK_W{delay_stage_select[112]}})
                                | (tmp_icb_cmd_pack_113 & {BUF_CMD_PACK_W{delay_stage_select[113]}})
                                | (tmp_icb_cmd_pack_114 & {BUF_CMD_PACK_W{delay_stage_select[114]}})
                                | (tmp_icb_cmd_pack_115 & {BUF_CMD_PACK_W{delay_stage_select[115]}})
                                | (tmp_icb_cmd_pack_116 & {BUF_CMD_PACK_W{delay_stage_select[116]}})
                                | (tmp_icb_cmd_pack_117 & {BUF_CMD_PACK_W{delay_stage_select[117]}})
                                | (tmp_icb_cmd_pack_118 & {BUF_CMD_PACK_W{delay_stage_select[118]}})
                                | (tmp_icb_cmd_pack_119 & {BUF_CMD_PACK_W{delay_stage_select[119]}})
                                | (tmp_icb_cmd_pack_120 & {BUF_CMD_PACK_W{delay_stage_select[120]}})
                                | (tmp_icb_cmd_pack_121 & {BUF_CMD_PACK_W{delay_stage_select[121]}})
                                | (tmp_icb_cmd_pack_122 & {BUF_CMD_PACK_W{delay_stage_select[122]}})
                                | (tmp_icb_cmd_pack_123 & {BUF_CMD_PACK_W{delay_stage_select[123]}})
                                | (tmp_icb_cmd_pack_124 & {BUF_CMD_PACK_W{delay_stage_select[124]}})
                                | (tmp_icb_cmd_pack_125 & {BUF_CMD_PACK_W{delay_stage_select[125]}})
                                | (tmp_icb_cmd_pack_126 & {BUF_CMD_PACK_W{delay_stage_select[126]}})
                                | (tmp_icb_cmd_pack_127 & {BUF_CMD_PACK_W{delay_stage_select[127]}})
                                | (tmp_icb_cmd_pack_128 & {BUF_CMD_PACK_W{delay_stage_select[128]}})
                                | (tmp_icb_cmd_pack_129 & {BUF_CMD_PACK_W{delay_stage_select[129]}})
                                | (tmp_icb_cmd_pack_130 & {BUF_CMD_PACK_W{delay_stage_select[130]}})
                                | (tmp_icb_cmd_pack_131 & {BUF_CMD_PACK_W{delay_stage_select[131]}})
                                | (tmp_icb_cmd_pack_132 & {BUF_CMD_PACK_W{delay_stage_select[132]}})
                                | (tmp_icb_cmd_pack_133 & {BUF_CMD_PACK_W{delay_stage_select[133]}})
                                | (tmp_icb_cmd_pack_134 & {BUF_CMD_PACK_W{delay_stage_select[134]}})
                                | (tmp_icb_cmd_pack_135 & {BUF_CMD_PACK_W{delay_stage_select[135]}})
                                | (tmp_icb_cmd_pack_136 & {BUF_CMD_PACK_W{delay_stage_select[136]}})
                                | (tmp_icb_cmd_pack_137 & {BUF_CMD_PACK_W{delay_stage_select[137]}})
                                | (tmp_icb_cmd_pack_138 & {BUF_CMD_PACK_W{delay_stage_select[138]}})
                                | (tmp_icb_cmd_pack_139 & {BUF_CMD_PACK_W{delay_stage_select[139]}})
                                | (tmp_icb_cmd_pack_140 & {BUF_CMD_PACK_W{delay_stage_select[140]}})
                                | (tmp_icb_cmd_pack_141 & {BUF_CMD_PACK_W{delay_stage_select[141]}})
                                | (tmp_icb_cmd_pack_142 & {BUF_CMD_PACK_W{delay_stage_select[142]}})
                                | (tmp_icb_cmd_pack_143 & {BUF_CMD_PACK_W{delay_stage_select[143]}})
                                | (tmp_icb_cmd_pack_144 & {BUF_CMD_PACK_W{delay_stage_select[144]}})
                                | (tmp_icb_cmd_pack_145 & {BUF_CMD_PACK_W{delay_stage_select[145]}})
                                | (tmp_icb_cmd_pack_146 & {BUF_CMD_PACK_W{delay_stage_select[146]}})
                                | (tmp_icb_cmd_pack_147 & {BUF_CMD_PACK_W{delay_stage_select[147]}})
                                | (tmp_icb_cmd_pack_148 & {BUF_CMD_PACK_W{delay_stage_select[148]}})
                                | (tmp_icb_cmd_pack_149 & {BUF_CMD_PACK_W{delay_stage_select[149]}})
                                | (tmp_icb_cmd_pack_150 & {BUF_CMD_PACK_W{delay_stage_select[150]}})
                                | (tmp_icb_cmd_pack_151 & {BUF_CMD_PACK_W{delay_stage_select[151]}})
                                | (tmp_icb_cmd_pack_152 & {BUF_CMD_PACK_W{delay_stage_select[152]}})
                                | (tmp_icb_cmd_pack_153 & {BUF_CMD_PACK_W{delay_stage_select[153]}})
                                | (tmp_icb_cmd_pack_154 & {BUF_CMD_PACK_W{delay_stage_select[154]}})
                                | (tmp_icb_cmd_pack_155 & {BUF_CMD_PACK_W{delay_stage_select[155]}})
                                | (tmp_icb_cmd_pack_156 & {BUF_CMD_PACK_W{delay_stage_select[156]}})
                                | (tmp_icb_cmd_pack_157 & {BUF_CMD_PACK_W{delay_stage_select[157]}})
                                | (tmp_icb_cmd_pack_158 & {BUF_CMD_PACK_W{delay_stage_select[158]}})
                                | (tmp_icb_cmd_pack_159 & {BUF_CMD_PACK_W{delay_stage_select[159]}})
                                | (tmp_icb_cmd_pack_160 & {BUF_CMD_PACK_W{delay_stage_select[160]}})
                                | (tmp_icb_cmd_pack_161 & {BUF_CMD_PACK_W{delay_stage_select[161]}})
                                | (tmp_icb_cmd_pack_162 & {BUF_CMD_PACK_W{delay_stage_select[162]}})
                                | (tmp_icb_cmd_pack_163 & {BUF_CMD_PACK_W{delay_stage_select[163]}})
                                | (tmp_icb_cmd_pack_164 & {BUF_CMD_PACK_W{delay_stage_select[164]}})
                                | (tmp_icb_cmd_pack_165 & {BUF_CMD_PACK_W{delay_stage_select[165]}})
                                | (tmp_icb_cmd_pack_166 & {BUF_CMD_PACK_W{delay_stage_select[166]}})
                                | (tmp_icb_cmd_pack_167 & {BUF_CMD_PACK_W{delay_stage_select[167]}})
                                | (tmp_icb_cmd_pack_168 & {BUF_CMD_PACK_W{delay_stage_select[168]}})
                                | (tmp_icb_cmd_pack_169 & {BUF_CMD_PACK_W{delay_stage_select[169]}})
                                | (tmp_icb_cmd_pack_170 & {BUF_CMD_PACK_W{delay_stage_select[170]}})
                                | (tmp_icb_cmd_pack_171 & {BUF_CMD_PACK_W{delay_stage_select[171]}})
                                | (tmp_icb_cmd_pack_172 & {BUF_CMD_PACK_W{delay_stage_select[172]}})
                                | (tmp_icb_cmd_pack_173 & {BUF_CMD_PACK_W{delay_stage_select[173]}})
                                | (tmp_icb_cmd_pack_174 & {BUF_CMD_PACK_W{delay_stage_select[174]}})
                                | (tmp_icb_cmd_pack_175 & {BUF_CMD_PACK_W{delay_stage_select[175]}})
                                | (tmp_icb_cmd_pack_176 & {BUF_CMD_PACK_W{delay_stage_select[176]}})
                                | (tmp_icb_cmd_pack_177 & {BUF_CMD_PACK_W{delay_stage_select[177]}})
                                | (tmp_icb_cmd_pack_178 & {BUF_CMD_PACK_W{delay_stage_select[178]}})
                                | (tmp_icb_cmd_pack_179 & {BUF_CMD_PACK_W{delay_stage_select[179]}})
                                | (tmp_icb_cmd_pack_180 & {BUF_CMD_PACK_W{delay_stage_select[180]}})
                                | (tmp_icb_cmd_pack_181 & {BUF_CMD_PACK_W{delay_stage_select[181]}})
                                | (tmp_icb_cmd_pack_182 & {BUF_CMD_PACK_W{delay_stage_select[182]}})
                                | (tmp_icb_cmd_pack_183 & {BUF_CMD_PACK_W{delay_stage_select[183]}})
                                | (tmp_icb_cmd_pack_184 & {BUF_CMD_PACK_W{delay_stage_select[184]}})
                                | (tmp_icb_cmd_pack_185 & {BUF_CMD_PACK_W{delay_stage_select[185]}})
                                | (tmp_icb_cmd_pack_186 & {BUF_CMD_PACK_W{delay_stage_select[186]}})
                                | (tmp_icb_cmd_pack_187 & {BUF_CMD_PACK_W{delay_stage_select[187]}})
                                | (tmp_icb_cmd_pack_188 & {BUF_CMD_PACK_W{delay_stage_select[188]}})
                                | (tmp_icb_cmd_pack_189 & {BUF_CMD_PACK_W{delay_stage_select[189]}})
                                | (tmp_icb_cmd_pack_190 & {BUF_CMD_PACK_W{delay_stage_select[190]}})
                                | (tmp_icb_cmd_pack_191 & {BUF_CMD_PACK_W{delay_stage_select[191]}})
                                | (tmp_icb_cmd_pack_192 & {BUF_CMD_PACK_W{delay_stage_select[192]}})
                                | (tmp_icb_cmd_pack_193 & {BUF_CMD_PACK_W{delay_stage_select[193]}})
                                | (tmp_icb_cmd_pack_194 & {BUF_CMD_PACK_W{delay_stage_select[194]}})
                                | (tmp_icb_cmd_pack_195 & {BUF_CMD_PACK_W{delay_stage_select[195]}})
                                | (tmp_icb_cmd_pack_196 & {BUF_CMD_PACK_W{delay_stage_select[196]}})
                                | (tmp_icb_cmd_pack_197 & {BUF_CMD_PACK_W{delay_stage_select[197]}})
                                | (tmp_icb_cmd_pack_198 & {BUF_CMD_PACK_W{delay_stage_select[198]}})
                                | (tmp_icb_cmd_pack_199 & {BUF_CMD_PACK_W{delay_stage_select[199]}})
                                | (tmp_icb_cmd_pack_200 & {BUF_CMD_PACK_W{delay_stage_select[200]}})
                                | (tmp_icb_cmd_pack_201 & {BUF_CMD_PACK_W{delay_stage_select[201]}})
                                | (tmp_icb_cmd_pack_202 & {BUF_CMD_PACK_W{delay_stage_select[202]}})
                                | (tmp_icb_cmd_pack_203 & {BUF_CMD_PACK_W{delay_stage_select[203]}})
                                | (tmp_icb_cmd_pack_204 & {BUF_CMD_PACK_W{delay_stage_select[204]}})
                                | (tmp_icb_cmd_pack_205 & {BUF_CMD_PACK_W{delay_stage_select[205]}})
                                | (tmp_icb_cmd_pack_206 & {BUF_CMD_PACK_W{delay_stage_select[206]}})
                                | (tmp_icb_cmd_pack_207 & {BUF_CMD_PACK_W{delay_stage_select[207]}})
                                | (tmp_icb_cmd_pack_208 & {BUF_CMD_PACK_W{delay_stage_select[208]}})
                                | (tmp_icb_cmd_pack_209 & {BUF_CMD_PACK_W{delay_stage_select[209]}})
                                | (tmp_icb_cmd_pack_210 & {BUF_CMD_PACK_W{delay_stage_select[210]}})
                                | (tmp_icb_cmd_pack_211 & {BUF_CMD_PACK_W{delay_stage_select[211]}})
                                | (tmp_icb_cmd_pack_212 & {BUF_CMD_PACK_W{delay_stage_select[212]}})
                                | (tmp_icb_cmd_pack_213 & {BUF_CMD_PACK_W{delay_stage_select[213]}})
                                | (tmp_icb_cmd_pack_214 & {BUF_CMD_PACK_W{delay_stage_select[214]}})
                                | (tmp_icb_cmd_pack_215 & {BUF_CMD_PACK_W{delay_stage_select[215]}})
                                | (tmp_icb_cmd_pack_216 & {BUF_CMD_PACK_W{delay_stage_select[216]}})
                                | (tmp_icb_cmd_pack_217 & {BUF_CMD_PACK_W{delay_stage_select[217]}})
                                | (tmp_icb_cmd_pack_218 & {BUF_CMD_PACK_W{delay_stage_select[218]}})
                                | (tmp_icb_cmd_pack_219 & {BUF_CMD_PACK_W{delay_stage_select[219]}})
                                | (tmp_icb_cmd_pack_220 & {BUF_CMD_PACK_W{delay_stage_select[220]}})
                                | (tmp_icb_cmd_pack_221 & {BUF_CMD_PACK_W{delay_stage_select[221]}})
                                | (tmp_icb_cmd_pack_222 & {BUF_CMD_PACK_W{delay_stage_select[222]}})
                                | (tmp_icb_cmd_pack_223 & {BUF_CMD_PACK_W{delay_stage_select[223]}})
                                | (tmp_icb_cmd_pack_224 & {BUF_CMD_PACK_W{delay_stage_select[224]}})
                                | (tmp_icb_cmd_pack_225 & {BUF_CMD_PACK_W{delay_stage_select[225]}})
                                | (tmp_icb_cmd_pack_226 & {BUF_CMD_PACK_W{delay_stage_select[226]}})
                                | (tmp_icb_cmd_pack_227 & {BUF_CMD_PACK_W{delay_stage_select[227]}})
                                | (tmp_icb_cmd_pack_228 & {BUF_CMD_PACK_W{delay_stage_select[228]}})
                                | (tmp_icb_cmd_pack_229 & {BUF_CMD_PACK_W{delay_stage_select[229]}})
                                | (tmp_icb_cmd_pack_230 & {BUF_CMD_PACK_W{delay_stage_select[230]}})
                                | (tmp_icb_cmd_pack_231 & {BUF_CMD_PACK_W{delay_stage_select[231]}})
                                | (tmp_icb_cmd_pack_232 & {BUF_CMD_PACK_W{delay_stage_select[232]}})
                                | (tmp_icb_cmd_pack_233 & {BUF_CMD_PACK_W{delay_stage_select[233]}})
                                | (tmp_icb_cmd_pack_234 & {BUF_CMD_PACK_W{delay_stage_select[234]}})
                                | (tmp_icb_cmd_pack_235 & {BUF_CMD_PACK_W{delay_stage_select[235]}})
                                | (tmp_icb_cmd_pack_236 & {BUF_CMD_PACK_W{delay_stage_select[236]}})
                                | (tmp_icb_cmd_pack_237 & {BUF_CMD_PACK_W{delay_stage_select[237]}})
                                | (tmp_icb_cmd_pack_238 & {BUF_CMD_PACK_W{delay_stage_select[238]}})
                                | (tmp_icb_cmd_pack_239 & {BUF_CMD_PACK_W{delay_stage_select[239]}})
                                | (tmp_icb_cmd_pack_240 & {BUF_CMD_PACK_W{delay_stage_select[240]}})
                                | (tmp_icb_cmd_pack_241 & {BUF_CMD_PACK_W{delay_stage_select[241]}})
                                | (tmp_icb_cmd_pack_242 & {BUF_CMD_PACK_W{delay_stage_select[242]}})
                                | (tmp_icb_cmd_pack_243 & {BUF_CMD_PACK_W{delay_stage_select[243]}})
                                | (tmp_icb_cmd_pack_244 & {BUF_CMD_PACK_W{delay_stage_select[244]}})
                                | (tmp_icb_cmd_pack_245 & {BUF_CMD_PACK_W{delay_stage_select[245]}})
                                | (tmp_icb_cmd_pack_246 & {BUF_CMD_PACK_W{delay_stage_select[246]}})
                                | (tmp_icb_cmd_pack_247 & {BUF_CMD_PACK_W{delay_stage_select[247]}})
                                | (tmp_icb_cmd_pack_248 & {BUF_CMD_PACK_W{delay_stage_select[248]}})
                                | (tmp_icb_cmd_pack_249 & {BUF_CMD_PACK_W{delay_stage_select[249]}})
                                | (tmp_icb_cmd_pack_250 & {BUF_CMD_PACK_W{delay_stage_select[250]}})
                                | (tmp_icb_cmd_pack_251 & {BUF_CMD_PACK_W{delay_stage_select[251]}})
                                | (tmp_icb_cmd_pack_252 & {BUF_CMD_PACK_W{delay_stage_select[252]}})
                                | (tmp_icb_cmd_pack_253 & {BUF_CMD_PACK_W{delay_stage_select[253]}})
                                | (tmp_icb_cmd_pack_254 & {BUF_CMD_PACK_W{delay_stage_select[254]}})
                                | (tmp_icb_cmd_pack_255 & {BUF_CMD_PACK_W{delay_stage_select[255]}})
                                | (tmp_icb_cmd_pack_256 & {BUF_CMD_PACK_W{delay_stage_select[256]}})
                                | (tmp_icb_cmd_pack_257 & {BUF_CMD_PACK_W{delay_stage_select[257]}})
                                | (tmp_icb_cmd_pack_258 & {BUF_CMD_PACK_W{delay_stage_select[258]}})
                                | (tmp_icb_cmd_pack_259 & {BUF_CMD_PACK_W{delay_stage_select[259]}})
                                | (tmp_icb_cmd_pack_260 & {BUF_CMD_PACK_W{delay_stage_select[260]}})
                                | (tmp_icb_cmd_pack_261 & {BUF_CMD_PACK_W{delay_stage_select[261]}})
                                | (tmp_icb_cmd_pack_262 & {BUF_CMD_PACK_W{delay_stage_select[262]}})
                                | (tmp_icb_cmd_pack_263 & {BUF_CMD_PACK_W{delay_stage_select[263]}})
                                | (tmp_icb_cmd_pack_264 & {BUF_CMD_PACK_W{delay_stage_select[264]}})
                                | (tmp_icb_cmd_pack_265 & {BUF_CMD_PACK_W{delay_stage_select[265]}})
                                | (tmp_icb_cmd_pack_266 & {BUF_CMD_PACK_W{delay_stage_select[266]}})
                                | (tmp_icb_cmd_pack_267 & {BUF_CMD_PACK_W{delay_stage_select[267]}})
                                | (tmp_icb_cmd_pack_268 & {BUF_CMD_PACK_W{delay_stage_select[268]}})
                                | (tmp_icb_cmd_pack_269 & {BUF_CMD_PACK_W{delay_stage_select[269]}})
                                | (tmp_icb_cmd_pack_270 & {BUF_CMD_PACK_W{delay_stage_select[270]}})
                                | (tmp_icb_cmd_pack_271 & {BUF_CMD_PACK_W{delay_stage_select[271]}})
                                | (tmp_icb_cmd_pack_272 & {BUF_CMD_PACK_W{delay_stage_select[272]}})
                                | (tmp_icb_cmd_pack_273 & {BUF_CMD_PACK_W{delay_stage_select[273]}})
                                | (tmp_icb_cmd_pack_274 & {BUF_CMD_PACK_W{delay_stage_select[274]}})
                                | (tmp_icb_cmd_pack_275 & {BUF_CMD_PACK_W{delay_stage_select[275]}})
                                | (tmp_icb_cmd_pack_276 & {BUF_CMD_PACK_W{delay_stage_select[276]}})
                                | (tmp_icb_cmd_pack_277 & {BUF_CMD_PACK_W{delay_stage_select[277]}})
                                | (tmp_icb_cmd_pack_278 & {BUF_CMD_PACK_W{delay_stage_select[278]}})
                                | (tmp_icb_cmd_pack_279 & {BUF_CMD_PACK_W{delay_stage_select[279]}})
                                | (tmp_icb_cmd_pack_280 & {BUF_CMD_PACK_W{delay_stage_select[280]}})
                                | (tmp_icb_cmd_pack_281 & {BUF_CMD_PACK_W{delay_stage_select[281]}})
                                | (tmp_icb_cmd_pack_282 & {BUF_CMD_PACK_W{delay_stage_select[282]}})
                                | (tmp_icb_cmd_pack_283 & {BUF_CMD_PACK_W{delay_stage_select[283]}})
                                | (tmp_icb_cmd_pack_284 & {BUF_CMD_PACK_W{delay_stage_select[284]}})
                                | (tmp_icb_cmd_pack_285 & {BUF_CMD_PACK_W{delay_stage_select[285]}})
                                | (tmp_icb_cmd_pack_286 & {BUF_CMD_PACK_W{delay_stage_select[286]}})
                                | (tmp_icb_cmd_pack_287 & {BUF_CMD_PACK_W{delay_stage_select[287]}})
                                | (tmp_icb_cmd_pack_288 & {BUF_CMD_PACK_W{delay_stage_select[288]}})
                                | (tmp_icb_cmd_pack_289 & {BUF_CMD_PACK_W{delay_stage_select[289]}})
                                | (tmp_icb_cmd_pack_290 & {BUF_CMD_PACK_W{delay_stage_select[290]}})
                                | (tmp_icb_cmd_pack_291 & {BUF_CMD_PACK_W{delay_stage_select[291]}})
                                | (tmp_icb_cmd_pack_292 & {BUF_CMD_PACK_W{delay_stage_select[292]}})
                                | (tmp_icb_cmd_pack_293 & {BUF_CMD_PACK_W{delay_stage_select[293]}})
                                | (tmp_icb_cmd_pack_294 & {BUF_CMD_PACK_W{delay_stage_select[294]}})
                                | (tmp_icb_cmd_pack_295 & {BUF_CMD_PACK_W{delay_stage_select[295]}})
                                | (tmp_icb_cmd_pack_296 & {BUF_CMD_PACK_W{delay_stage_select[296]}})
                                | (tmp_icb_cmd_pack_297 & {BUF_CMD_PACK_W{delay_stage_select[297]}})
                                | (tmp_icb_cmd_pack_298 & {BUF_CMD_PACK_W{delay_stage_select[298]}})
                                | (tmp_icb_cmd_pack_299 & {BUF_CMD_PACK_W{delay_stage_select[299]}})
                                | (tmp_icb_cmd_pack_300 & {BUF_CMD_PACK_W{delay_stage_select[300]}})
                                | (tmp_icb_cmd_pack_301 & {BUF_CMD_PACK_W{delay_stage_select[301]}})
                                | (tmp_icb_cmd_pack_302 & {BUF_CMD_PACK_W{delay_stage_select[302]}})
                                | (tmp_icb_cmd_pack_303 & {BUF_CMD_PACK_W{delay_stage_select[303]}})
                                | (tmp_icb_cmd_pack_304 & {BUF_CMD_PACK_W{delay_stage_select[304]}})
                                | (tmp_icb_cmd_pack_305 & {BUF_CMD_PACK_W{delay_stage_select[305]}})
                                | (tmp_icb_cmd_pack_306 & {BUF_CMD_PACK_W{delay_stage_select[306]}})
                                | (tmp_icb_cmd_pack_307 & {BUF_CMD_PACK_W{delay_stage_select[307]}})
                                | (tmp_icb_cmd_pack_308 & {BUF_CMD_PACK_W{delay_stage_select[308]}})
                                | (tmp_icb_cmd_pack_309 & {BUF_CMD_PACK_W{delay_stage_select[309]}})
                                | (tmp_icb_cmd_pack_310 & {BUF_CMD_PACK_W{delay_stage_select[310]}})
                                | (tmp_icb_cmd_pack_311 & {BUF_CMD_PACK_W{delay_stage_select[311]}})
                                | (tmp_icb_cmd_pack_312 & {BUF_CMD_PACK_W{delay_stage_select[312]}})
                                | (tmp_icb_cmd_pack_313 & {BUF_CMD_PACK_W{delay_stage_select[313]}})
                                | (tmp_icb_cmd_pack_314 & {BUF_CMD_PACK_W{delay_stage_select[314]}})
                                | (tmp_icb_cmd_pack_315 & {BUF_CMD_PACK_W{delay_stage_select[315]}})
                                | (tmp_icb_cmd_pack_316 & {BUF_CMD_PACK_W{delay_stage_select[316]}})
                                | (tmp_icb_cmd_pack_317 & {BUF_CMD_PACK_W{delay_stage_select[317]}})
                                | (tmp_icb_cmd_pack_318 & {BUF_CMD_PACK_W{delay_stage_select[318]}})
                                | (tmp_icb_cmd_pack_319 & {BUF_CMD_PACK_W{delay_stage_select[319]}})
                                | (tmp_icb_cmd_pack_320 & {BUF_CMD_PACK_W{delay_stage_select[320]}})
                                | (tmp_icb_cmd_pack_321 & {BUF_CMD_PACK_W{delay_stage_select[321]}})
                                | (tmp_icb_cmd_pack_322 & {BUF_CMD_PACK_W{delay_stage_select[322]}})
                                | (tmp_icb_cmd_pack_323 & {BUF_CMD_PACK_W{delay_stage_select[323]}})
                                | (tmp_icb_cmd_pack_324 & {BUF_CMD_PACK_W{delay_stage_select[324]}})
                                | (tmp_icb_cmd_pack_325 & {BUF_CMD_PACK_W{delay_stage_select[325]}})
                                | (tmp_icb_cmd_pack_326 & {BUF_CMD_PACK_W{delay_stage_select[326]}})
                                | (tmp_icb_cmd_pack_327 & {BUF_CMD_PACK_W{delay_stage_select[327]}})
                                | (tmp_icb_cmd_pack_328 & {BUF_CMD_PACK_W{delay_stage_select[328]}})
                                | (tmp_icb_cmd_pack_329 & {BUF_CMD_PACK_W{delay_stage_select[329]}})
                                | (tmp_icb_cmd_pack_330 & {BUF_CMD_PACK_W{delay_stage_select[330]}})
                                | (tmp_icb_cmd_pack_331 & {BUF_CMD_PACK_W{delay_stage_select[331]}})
                                | (tmp_icb_cmd_pack_332 & {BUF_CMD_PACK_W{delay_stage_select[332]}})
                                | (tmp_icb_cmd_pack_333 & {BUF_CMD_PACK_W{delay_stage_select[333]}})
                                | (tmp_icb_cmd_pack_334 & {BUF_CMD_PACK_W{delay_stage_select[334]}})
                                | (tmp_icb_cmd_pack_335 & {BUF_CMD_PACK_W{delay_stage_select[335]}})
                                | (tmp_icb_cmd_pack_336 & {BUF_CMD_PACK_W{delay_stage_select[336]}})
                                | (tmp_icb_cmd_pack_337 & {BUF_CMD_PACK_W{delay_stage_select[337]}})
                                | (tmp_icb_cmd_pack_338 & {BUF_CMD_PACK_W{delay_stage_select[338]}})
                                | (tmp_icb_cmd_pack_339 & {BUF_CMD_PACK_W{delay_stage_select[339]}})
                                | (tmp_icb_cmd_pack_340 & {BUF_CMD_PACK_W{delay_stage_select[340]}})
                                | (tmp_icb_cmd_pack_341 & {BUF_CMD_PACK_W{delay_stage_select[341]}})
                                | (tmp_icb_cmd_pack_342 & {BUF_CMD_PACK_W{delay_stage_select[342]}})
                                | (tmp_icb_cmd_pack_343 & {BUF_CMD_PACK_W{delay_stage_select[343]}})
                                | (tmp_icb_cmd_pack_344 & {BUF_CMD_PACK_W{delay_stage_select[344]}})
                                | (tmp_icb_cmd_pack_345 & {BUF_CMD_PACK_W{delay_stage_select[345]}})
                                | (tmp_icb_cmd_pack_346 & {BUF_CMD_PACK_W{delay_stage_select[346]}})
                                | (tmp_icb_cmd_pack_347 & {BUF_CMD_PACK_W{delay_stage_select[347]}})
                                | (tmp_icb_cmd_pack_348 & {BUF_CMD_PACK_W{delay_stage_select[348]}})
                                | (tmp_icb_cmd_pack_349 & {BUF_CMD_PACK_W{delay_stage_select[349]}})
                                | (tmp_icb_cmd_pack_350 & {BUF_CMD_PACK_W{delay_stage_select[350]}})
                                | (tmp_icb_cmd_pack_351 & {BUF_CMD_PACK_W{delay_stage_select[351]}})
                                | (tmp_icb_cmd_pack_352 & {BUF_CMD_PACK_W{delay_stage_select[352]}})
                                | (tmp_icb_cmd_pack_353 & {BUF_CMD_PACK_W{delay_stage_select[353]}})
                                | (tmp_icb_cmd_pack_354 & {BUF_CMD_PACK_W{delay_stage_select[354]}})
                                | (tmp_icb_cmd_pack_355 & {BUF_CMD_PACK_W{delay_stage_select[355]}})
                                | (tmp_icb_cmd_pack_356 & {BUF_CMD_PACK_W{delay_stage_select[356]}})
                                | (tmp_icb_cmd_pack_357 & {BUF_CMD_PACK_W{delay_stage_select[357]}})
                                | (tmp_icb_cmd_pack_358 & {BUF_CMD_PACK_W{delay_stage_select[358]}})
                                | (tmp_icb_cmd_pack_359 & {BUF_CMD_PACK_W{delay_stage_select[359]}})
                                | (tmp_icb_cmd_pack_360 & {BUF_CMD_PACK_W{delay_stage_select[360]}})
                                | (tmp_icb_cmd_pack_361 & {BUF_CMD_PACK_W{delay_stage_select[361]}})
                                | (tmp_icb_cmd_pack_362 & {BUF_CMD_PACK_W{delay_stage_select[362]}})
                                | (tmp_icb_cmd_pack_363 & {BUF_CMD_PACK_W{delay_stage_select[363]}})
                                | (tmp_icb_cmd_pack_364 & {BUF_CMD_PACK_W{delay_stage_select[364]}})
                                | (tmp_icb_cmd_pack_365 & {BUF_CMD_PACK_W{delay_stage_select[365]}})
                                | (tmp_icb_cmd_pack_366 & {BUF_CMD_PACK_W{delay_stage_select[366]}})
                                | (tmp_icb_cmd_pack_367 & {BUF_CMD_PACK_W{delay_stage_select[367]}})
                                | (tmp_icb_cmd_pack_368 & {BUF_CMD_PACK_W{delay_stage_select[368]}})
                                | (tmp_icb_cmd_pack_369 & {BUF_CMD_PACK_W{delay_stage_select[369]}})
                                | (tmp_icb_cmd_pack_370 & {BUF_CMD_PACK_W{delay_stage_select[370]}})
                                | (tmp_icb_cmd_pack_371 & {BUF_CMD_PACK_W{delay_stage_select[371]}})
                                | (tmp_icb_cmd_pack_372 & {BUF_CMD_PACK_W{delay_stage_select[372]}})
                                | (tmp_icb_cmd_pack_373 & {BUF_CMD_PACK_W{delay_stage_select[373]}})
                                | (tmp_icb_cmd_pack_374 & {BUF_CMD_PACK_W{delay_stage_select[374]}})
                                | (tmp_icb_cmd_pack_375 & {BUF_CMD_PACK_W{delay_stage_select[375]}})
                                | (tmp_icb_cmd_pack_376 & {BUF_CMD_PACK_W{delay_stage_select[376]}})
                                | (tmp_icb_cmd_pack_377 & {BUF_CMD_PACK_W{delay_stage_select[377]}})
                                | (tmp_icb_cmd_pack_378 & {BUF_CMD_PACK_W{delay_stage_select[378]}})
                                | (tmp_icb_cmd_pack_379 & {BUF_CMD_PACK_W{delay_stage_select[379]}})
                                | (tmp_icb_cmd_pack_380 & {BUF_CMD_PACK_W{delay_stage_select[380]}})
                                | (tmp_icb_cmd_pack_381 & {BUF_CMD_PACK_W{delay_stage_select[381]}})
                                | (tmp_icb_cmd_pack_382 & {BUF_CMD_PACK_W{delay_stage_select[382]}})
                                | (tmp_icb_cmd_pack_383 & {BUF_CMD_PACK_W{delay_stage_select[383]}})
                                | (tmp_icb_cmd_pack_384 & {BUF_CMD_PACK_W{delay_stage_select[384]}})
                                | (tmp_icb_cmd_pack_385 & {BUF_CMD_PACK_W{delay_stage_select[385]}})
                                | (tmp_icb_cmd_pack_386 & {BUF_CMD_PACK_W{delay_stage_select[386]}})
                                | (tmp_icb_cmd_pack_387 & {BUF_CMD_PACK_W{delay_stage_select[387]}})
                                | (tmp_icb_cmd_pack_388 & {BUF_CMD_PACK_W{delay_stage_select[388]}})
                                | (tmp_icb_cmd_pack_389 & {BUF_CMD_PACK_W{delay_stage_select[389]}})
                                | (tmp_icb_cmd_pack_390 & {BUF_CMD_PACK_W{delay_stage_select[390]}})
                                | (tmp_icb_cmd_pack_391 & {BUF_CMD_PACK_W{delay_stage_select[391]}})
                                | (tmp_icb_cmd_pack_392 & {BUF_CMD_PACK_W{delay_stage_select[392]}})
                                | (tmp_icb_cmd_pack_393 & {BUF_CMD_PACK_W{delay_stage_select[393]}})
                                | (tmp_icb_cmd_pack_394 & {BUF_CMD_PACK_W{delay_stage_select[394]}})
                                | (tmp_icb_cmd_pack_395 & {BUF_CMD_PACK_W{delay_stage_select[395]}})
                                | (tmp_icb_cmd_pack_396 & {BUF_CMD_PACK_W{delay_stage_select[396]}})
                                | (tmp_icb_cmd_pack_397 & {BUF_CMD_PACK_W{delay_stage_select[397]}})
                                | (tmp_icb_cmd_pack_398 & {BUF_CMD_PACK_W{delay_stage_select[398]}})
                                | (tmp_icb_cmd_pack_399 & {BUF_CMD_PACK_W{delay_stage_select[399]}})
                                | (tmp_icb_cmd_pack_400 & {BUF_CMD_PACK_W{delay_stage_select[400]}})
                                | (tmp_icb_cmd_pack_401 & {BUF_CMD_PACK_W{delay_stage_select[401]}})
                                | (tmp_icb_cmd_pack_402 & {BUF_CMD_PACK_W{delay_stage_select[402]}})
                                | (tmp_icb_cmd_pack_403 & {BUF_CMD_PACK_W{delay_stage_select[403]}})
                                | (tmp_icb_cmd_pack_404 & {BUF_CMD_PACK_W{delay_stage_select[404]}})
                                | (tmp_icb_cmd_pack_405 & {BUF_CMD_PACK_W{delay_stage_select[405]}})
                                | (tmp_icb_cmd_pack_406 & {BUF_CMD_PACK_W{delay_stage_select[406]}})
                                | (tmp_icb_cmd_pack_407 & {BUF_CMD_PACK_W{delay_stage_select[407]}})
                                | (tmp_icb_cmd_pack_408 & {BUF_CMD_PACK_W{delay_stage_select[408]}})
                                | (tmp_icb_cmd_pack_409 & {BUF_CMD_PACK_W{delay_stage_select[409]}})
                                | (tmp_icb_cmd_pack_410 & {BUF_CMD_PACK_W{delay_stage_select[410]}})
                                | (tmp_icb_cmd_pack_411 & {BUF_CMD_PACK_W{delay_stage_select[411]}})
                                | (tmp_icb_cmd_pack_412 & {BUF_CMD_PACK_W{delay_stage_select[412]}})
                                | (tmp_icb_cmd_pack_413 & {BUF_CMD_PACK_W{delay_stage_select[413]}})
                                | (tmp_icb_cmd_pack_414 & {BUF_CMD_PACK_W{delay_stage_select[414]}})
                                | (tmp_icb_cmd_pack_415 & {BUF_CMD_PACK_W{delay_stage_select[415]}})
                                | (tmp_icb_cmd_pack_416 & {BUF_CMD_PACK_W{delay_stage_select[416]}})
                                | (tmp_icb_cmd_pack_417 & {BUF_CMD_PACK_W{delay_stage_select[417]}})
                                | (tmp_icb_cmd_pack_418 & {BUF_CMD_PACK_W{delay_stage_select[418]}})
                                | (tmp_icb_cmd_pack_419 & {BUF_CMD_PACK_W{delay_stage_select[419]}})
                                | (tmp_icb_cmd_pack_420 & {BUF_CMD_PACK_W{delay_stage_select[420]}})
                                | (tmp_icb_cmd_pack_421 & {BUF_CMD_PACK_W{delay_stage_select[421]}})
                                | (tmp_icb_cmd_pack_422 & {BUF_CMD_PACK_W{delay_stage_select[422]}})
                                | (tmp_icb_cmd_pack_423 & {BUF_CMD_PACK_W{delay_stage_select[423]}})
                                | (tmp_icb_cmd_pack_424 & {BUF_CMD_PACK_W{delay_stage_select[424]}})
                                | (tmp_icb_cmd_pack_425 & {BUF_CMD_PACK_W{delay_stage_select[425]}})
                                | (tmp_icb_cmd_pack_426 & {BUF_CMD_PACK_W{delay_stage_select[426]}})
                                | (tmp_icb_cmd_pack_427 & {BUF_CMD_PACK_W{delay_stage_select[427]}})
                                | (tmp_icb_cmd_pack_428 & {BUF_CMD_PACK_W{delay_stage_select[428]}})
                                | (tmp_icb_cmd_pack_429 & {BUF_CMD_PACK_W{delay_stage_select[429]}})
                                | (tmp_icb_cmd_pack_430 & {BUF_CMD_PACK_W{delay_stage_select[430]}})
                                | (tmp_icb_cmd_pack_431 & {BUF_CMD_PACK_W{delay_stage_select[431]}})
                                | (tmp_icb_cmd_pack_432 & {BUF_CMD_PACK_W{delay_stage_select[432]}})
                                | (tmp_icb_cmd_pack_433 & {BUF_CMD_PACK_W{delay_stage_select[433]}})
                                | (tmp_icb_cmd_pack_434 & {BUF_CMD_PACK_W{delay_stage_select[434]}})
                                | (tmp_icb_cmd_pack_435 & {BUF_CMD_PACK_W{delay_stage_select[435]}})
                                | (tmp_icb_cmd_pack_436 & {BUF_CMD_PACK_W{delay_stage_select[436]}})
                                | (tmp_icb_cmd_pack_437 & {BUF_CMD_PACK_W{delay_stage_select[437]}})
                                | (tmp_icb_cmd_pack_438 & {BUF_CMD_PACK_W{delay_stage_select[438]}})
                                | (tmp_icb_cmd_pack_439 & {BUF_CMD_PACK_W{delay_stage_select[439]}})
                                | (tmp_icb_cmd_pack_440 & {BUF_CMD_PACK_W{delay_stage_select[440]}})
                                | (tmp_icb_cmd_pack_441 & {BUF_CMD_PACK_W{delay_stage_select[441]}})
                                | (tmp_icb_cmd_pack_442 & {BUF_CMD_PACK_W{delay_stage_select[442]}})
                                | (tmp_icb_cmd_pack_443 & {BUF_CMD_PACK_W{delay_stage_select[443]}})
                                | (tmp_icb_cmd_pack_444 & {BUF_CMD_PACK_W{delay_stage_select[444]}})
                                | (tmp_icb_cmd_pack_445 & {BUF_CMD_PACK_W{delay_stage_select[445]}})
                                | (tmp_icb_cmd_pack_446 & {BUF_CMD_PACK_W{delay_stage_select[446]}})
                                | (tmp_icb_cmd_pack_447 & {BUF_CMD_PACK_W{delay_stage_select[447]}})
                                | (tmp_icb_cmd_pack_448 & {BUF_CMD_PACK_W{delay_stage_select[448]}})
                                | (tmp_icb_cmd_pack_449 & {BUF_CMD_PACK_W{delay_stage_select[449]}})
                                | (tmp_icb_cmd_pack_450 & {BUF_CMD_PACK_W{delay_stage_select[450]}})
                                | (tmp_icb_cmd_pack_451 & {BUF_CMD_PACK_W{delay_stage_select[451]}})
                                | (tmp_icb_cmd_pack_452 & {BUF_CMD_PACK_W{delay_stage_select[452]}})
                                | (tmp_icb_cmd_pack_453 & {BUF_CMD_PACK_W{delay_stage_select[453]}})
                                | (tmp_icb_cmd_pack_454 & {BUF_CMD_PACK_W{delay_stage_select[454]}})
                                | (tmp_icb_cmd_pack_455 & {BUF_CMD_PACK_W{delay_stage_select[455]}})
                                | (tmp_icb_cmd_pack_456 & {BUF_CMD_PACK_W{delay_stage_select[456]}})
                                | (tmp_icb_cmd_pack_457 & {BUF_CMD_PACK_W{delay_stage_select[457]}})
                                | (tmp_icb_cmd_pack_458 & {BUF_CMD_PACK_W{delay_stage_select[458]}})
                                | (tmp_icb_cmd_pack_459 & {BUF_CMD_PACK_W{delay_stage_select[459]}})
                                | (tmp_icb_cmd_pack_460 & {BUF_CMD_PACK_W{delay_stage_select[460]}})
                                | (tmp_icb_cmd_pack_461 & {BUF_CMD_PACK_W{delay_stage_select[461]}})
                                | (tmp_icb_cmd_pack_462 & {BUF_CMD_PACK_W{delay_stage_select[462]}})
                                | (tmp_icb_cmd_pack_463 & {BUF_CMD_PACK_W{delay_stage_select[463]}})
                                | (tmp_icb_cmd_pack_464 & {BUF_CMD_PACK_W{delay_stage_select[464]}})
                                | (tmp_icb_cmd_pack_465 & {BUF_CMD_PACK_W{delay_stage_select[465]}})
                                | (tmp_icb_cmd_pack_466 & {BUF_CMD_PACK_W{delay_stage_select[466]}})
                                | (tmp_icb_cmd_pack_467 & {BUF_CMD_PACK_W{delay_stage_select[467]}})
                                | (tmp_icb_cmd_pack_468 & {BUF_CMD_PACK_W{delay_stage_select[468]}})
                                | (tmp_icb_cmd_pack_469 & {BUF_CMD_PACK_W{delay_stage_select[469]}})
                                | (tmp_icb_cmd_pack_470 & {BUF_CMD_PACK_W{delay_stage_select[470]}})
                                | (tmp_icb_cmd_pack_471 & {BUF_CMD_PACK_W{delay_stage_select[471]}})
                                | (tmp_icb_cmd_pack_472 & {BUF_CMD_PACK_W{delay_stage_select[472]}})
                                | (tmp_icb_cmd_pack_473 & {BUF_CMD_PACK_W{delay_stage_select[473]}})
                                | (tmp_icb_cmd_pack_474 & {BUF_CMD_PACK_W{delay_stage_select[474]}})
                                | (tmp_icb_cmd_pack_475 & {BUF_CMD_PACK_W{delay_stage_select[475]}})
                                | (tmp_icb_cmd_pack_476 & {BUF_CMD_PACK_W{delay_stage_select[476]}})
                                | (tmp_icb_cmd_pack_477 & {BUF_CMD_PACK_W{delay_stage_select[477]}})
                                | (tmp_icb_cmd_pack_478 & {BUF_CMD_PACK_W{delay_stage_select[478]}})
                                | (tmp_icb_cmd_pack_479 & {BUF_CMD_PACK_W{delay_stage_select[479]}})
                                | (tmp_icb_cmd_pack_480 & {BUF_CMD_PACK_W{delay_stage_select[480]}})
                                | (tmp_icb_cmd_pack_481 & {BUF_CMD_PACK_W{delay_stage_select[481]}})
                                | (tmp_icb_cmd_pack_482 & {BUF_CMD_PACK_W{delay_stage_select[482]}})
                                | (tmp_icb_cmd_pack_483 & {BUF_CMD_PACK_W{delay_stage_select[483]}})
                                | (tmp_icb_cmd_pack_484 & {BUF_CMD_PACK_W{delay_stage_select[484]}})
                                | (tmp_icb_cmd_pack_485 & {BUF_CMD_PACK_W{delay_stage_select[485]}})
                                | (tmp_icb_cmd_pack_486 & {BUF_CMD_PACK_W{delay_stage_select[486]}})
                                | (tmp_icb_cmd_pack_487 & {BUF_CMD_PACK_W{delay_stage_select[487]}})
                                | (tmp_icb_cmd_pack_488 & {BUF_CMD_PACK_W{delay_stage_select[488]}})
                                | (tmp_icb_cmd_pack_489 & {BUF_CMD_PACK_W{delay_stage_select[489]}})
                                | (tmp_icb_cmd_pack_490 & {BUF_CMD_PACK_W{delay_stage_select[490]}})
                                | (tmp_icb_cmd_pack_491 & {BUF_CMD_PACK_W{delay_stage_select[491]}})
                                | (tmp_icb_cmd_pack_492 & {BUF_CMD_PACK_W{delay_stage_select[492]}})
                                | (tmp_icb_cmd_pack_493 & {BUF_CMD_PACK_W{delay_stage_select[493]}})
                                | (tmp_icb_cmd_pack_494 & {BUF_CMD_PACK_W{delay_stage_select[494]}})
                                | (tmp_icb_cmd_pack_495 & {BUF_CMD_PACK_W{delay_stage_select[495]}})
                                | (tmp_icb_cmd_pack_496 & {BUF_CMD_PACK_W{delay_stage_select[496]}})
                                | (tmp_icb_cmd_pack_497 & {BUF_CMD_PACK_W{delay_stage_select[497]}})
                                | (tmp_icb_cmd_pack_498 & {BUF_CMD_PACK_W{delay_stage_select[498]}})
                                | (tmp_icb_cmd_pack_499 & {BUF_CMD_PACK_W{delay_stage_select[499]}})
                                | (tmp_icb_cmd_pack_500 & {BUF_CMD_PACK_W{delay_stage_select[500]}})
                                | (tmp_icb_cmd_pack_501 & {BUF_CMD_PACK_W{delay_stage_select[501]}})
                                | (tmp_icb_cmd_pack_502 & {BUF_CMD_PACK_W{delay_stage_select[502]}})
                                | (tmp_icb_cmd_pack_503 & {BUF_CMD_PACK_W{delay_stage_select[503]}})
                                | (tmp_icb_cmd_pack_504 & {BUF_CMD_PACK_W{delay_stage_select[504]}})
                                | (tmp_icb_cmd_pack_505 & {BUF_CMD_PACK_W{delay_stage_select[505]}})
                                | (tmp_icb_cmd_pack_506 & {BUF_CMD_PACK_W{delay_stage_select[506]}})
                                | (tmp_icb_cmd_pack_507 & {BUF_CMD_PACK_W{delay_stage_select[507]}})
                                | (tmp_icb_cmd_pack_508 & {BUF_CMD_PACK_W{delay_stage_select[508]}})
                                | (tmp_icb_cmd_pack_509 & {BUF_CMD_PACK_W{delay_stage_select[509]}})
                                | (tmp_icb_cmd_pack_510 & {BUF_CMD_PACK_W{delay_stage_select[510]}})
                                | (tmp_icb_cmd_pack_511 & {BUF_CMD_PACK_W{delay_stage_select[511]}})
                                ;
`endif
`endif 
  assign o_icb_cmd_valid    = byp_icb_cmd_valid; 
  assign byp_icb_cmd_ready  = o_icb_cmd_ready; 
  assign o_icb_cmd_read     = byp_icb_cmd_read; 
  assign o_icb_cmd_addr     = byp_icb_cmd_addr;  
  assign o_icb_cmd_wdata    = byp_icb_cmd_wdata; 
  assign o_icb_cmd_wmask    = byp_icb_cmd_wmask; 
  assign o_icb_cmd_usr      = byp_icb_cmd_usr;   
endmodule
