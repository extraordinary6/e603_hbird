 /*                                                                      
  *  Copyright (c) 2018-2025 Nuclei System Technology, Inc.       
  *  All rights reserved.                                                
  */                                                                     
module e603_subsys_bus_fab (
  input              i_axi_arvalid                 ,
  output             i_axi_arready                 ,
  input  [  31:   0] i_axi_araddr                  ,
  input  [   7:   0] i_axi_arlen                   ,
  input  [   2:   0] i_axi_arsize                  ,
  input  [   1:   0] i_axi_arburst                 ,
  input              i_axi_arlock                  ,
  input  [   3:   0] i_axi_arcache                 ,
  input  [   2:   0] i_axi_arprot                  ,
  input              i_axi_rready                  ,
  output             i_axi_rvalid                  ,
  output [  63:   0] i_axi_rdata                   ,
  output [   1:   0] i_axi_rresp                   ,
  output             i_axi_rlast                   ,
  input              i_axi_awvalid                 ,
  output             i_axi_awready                 ,
  input  [  31:   0] i_axi_awaddr                  ,
  input  [   7:   0] i_axi_awlen                   ,
  input  [   2:   0] i_axi_awsize                  ,
  input  [   1:   0] i_axi_awburst                 ,
  input              i_axi_awlock                  ,
  input  [   3:   0] i_axi_awcache                 ,
  input  [   2:   0] i_axi_awprot                  ,
  input              i_axi_bready                  ,
  output             i_axi_bvalid                  ,
  output [   1:   0] i_axi_bresp                   ,
  output             i_axi_wready                  ,
  input              i_axi_wvalid                  ,
  input  [  63:   0] i_axi_wdata                   ,
  input  [   7:   0] i_axi_wstrb                   ,
  input              i_axi_wlast                   ,
  input              udma_r_icb_cmd_valid          ,
  output             udma_r_icb_cmd_ready          ,
  input              udma_r_icb_cmd_sel            ,
  input              udma_r_icb_cmd_read           ,
  input  [  31:   0] udma_r_icb_cmd_addr           ,
  input  [  63:   0] udma_r_icb_cmd_wdata          ,
  input  [   7:   0] udma_r_icb_cmd_wmask          ,
  input  [   2:   0] udma_r_icb_cmd_size           ,
  input              udma_r_icb_cmd_lock           ,
  input              udma_r_icb_cmd_excl           ,
  input  [   7:   0] udma_r_icb_cmd_xlen           ,
  input  [   1:   0] udma_r_icb_cmd_xburst         ,
  input  [   1:   0] udma_r_icb_cmd_modes          ,
  input              udma_r_icb_cmd_dmode          ,
  input  [   2:   0] udma_r_icb_cmd_attri          ,
  input  [   1:   0] udma_r_icb_cmd_beat           ,
  input              udma_r_icb_rsp_ready          ,
  output             udma_r_icb_rsp_valid          ,
  output             udma_r_icb_rsp_err            ,
  output             udma_r_icb_rsp_excl_ok        ,
  output [  63:   0] udma_r_icb_rsp_rdata          ,
  input              udma_w_icb_cmd_valid          ,
  output             udma_w_icb_cmd_ready          ,
  input              udma_w_icb_cmd_sel            ,
  input              udma_w_icb_cmd_read           ,
  input  [  31:   0] udma_w_icb_cmd_addr           ,
  input  [  63:   0] udma_w_icb_cmd_wdata          ,
  input  [   7:   0] udma_w_icb_cmd_wmask          ,
  input  [   2:   0] udma_w_icb_cmd_size           ,
  input              udma_w_icb_cmd_lock           ,
  input              udma_w_icb_cmd_excl           ,
  input  [   7:   0] udma_w_icb_cmd_xlen           ,
  input  [   1:   0] udma_w_icb_cmd_xburst         ,
  input  [   1:   0] udma_w_icb_cmd_modes          ,
  input              udma_w_icb_cmd_dmode          ,
  input  [   2:   0] udma_w_icb_cmd_attri          ,
  input  [   1:   0] udma_w_icb_cmd_beat           ,
  input              udma_w_icb_rsp_ready          ,
  output             udma_w_icb_rsp_valid          ,
  output             udma_w_icb_rsp_err            ,
  output             udma_w_icb_rsp_excl_ok        ,
  output [  63:   0] udma_w_icb_rsp_rdata          ,
  input              dummy_icb_cmd_valid           ,
  output             dummy_icb_cmd_ready           ,
  input              dummy_icb_cmd_sel             ,
  input              dummy_icb_cmd_read            ,
  input  [  31:   0] dummy_icb_cmd_addr            ,
  input  [  63:   0] dummy_icb_cmd_wdata           ,
  input  [   7:   0] dummy_icb_cmd_wmask           ,
  input  [   2:   0] dummy_icb_cmd_size            ,
  input              dummy_icb_cmd_lock            ,
  input              dummy_icb_cmd_excl            ,
  input  [   7:   0] dummy_icb_cmd_xlen            ,
  input  [   1:   0] dummy_icb_cmd_xburst          ,
  input  [   1:   0] dummy_icb_cmd_modes           ,
  input              dummy_icb_cmd_dmode           ,
  input  [   2:   0] dummy_icb_cmd_attri           ,
  input  [   1:   0] dummy_icb_cmd_beat            ,
  input              dummy_icb_rsp_ready           ,
  output             dummy_icb_rsp_valid           ,
  output             dummy_icb_rsp_err             ,
  output             dummy_icb_rsp_excl_ok         ,
  output [  63:   0] dummy_icb_rsp_rdata           ,
  input              dummy_axi_arvalid             ,
  output             dummy_axi_arready             ,
  input  [  31:   0] dummy_axi_araddr              ,
  input  [   7:   0] dummy_axi_arlen               ,
  input  [   2:   0] dummy_axi_arsize              ,
  input  [   1:   0] dummy_axi_arburst             ,
  input              dummy_axi_arlock              ,
  input  [   3:   0] dummy_axi_arcache             ,
  input  [   2:   0] dummy_axi_arprot              ,
  input              dummy_axi_rready              ,
  output             dummy_axi_rvalid              ,
  output [  63:   0] dummy_axi_rdata               ,
  output [   1:   0] dummy_axi_rresp               ,
  output             dummy_axi_rlast               ,
  input              dummy_axi_awvalid             ,
  output             dummy_axi_awready             ,
  input  [  31:   0] dummy_axi_awaddr              ,
  input  [   7:   0] dummy_axi_awlen               ,
  input  [   2:   0] dummy_axi_awsize              ,
  input  [   1:   0] dummy_axi_awburst             ,
  input              dummy_axi_awlock              ,
  input  [   3:   0] dummy_axi_awcache             ,
  input  [   2:   0] dummy_axi_awprot              ,
  input              dummy_axi_bready              ,
  output             dummy_axi_bvalid              ,
  output [   1:   0] dummy_axi_bresp               ,
  output             dummy_axi_wready              ,
  input              dummy_axi_wvalid              ,
  input  [  63:   0] dummy_axi_wdata               ,
  input  [   7:   0] dummy_axi_wstrb               ,
  input              dummy_axi_wlast               ,
  input  [   1:   0] dummy_ahbl_htrans             ,
  input              dummy_ahbl_hwrite             ,
  input              dummy_ahbl_hmastlock          ,
  input  [   2:   0] dummy_ahbl_hsize              ,
  input  [   2:   0] dummy_ahbl_hburst             ,
  input  [   3:   0] dummy_ahbl_hprot              ,
  input  [  63:   0] dummy_ahbl_hwdata             ,
  input  [  31:   0] dummy_ahbl_haddr              ,
  output [  63:   0] dummy_ahbl_hrdata             ,
  output [   1:   0] dummy_ahbl_hresp              ,
  output             dummy_ahbl_hready             ,
  input              eth_axi_arvalid               ,
  output             eth_axi_arready               ,
  input  [  31:   0] eth_axi_araddr                ,
  input  [   7:   0] eth_axi_arlen                 ,
  input  [   2:   0] eth_axi_arsize                ,
  input  [   1:   0] eth_axi_arburst               ,
  input              eth_axi_arlock                ,
  input  [   3:   0] eth_axi_arcache               ,
  input  [   2:   0] eth_axi_arprot                ,
  input              eth_axi_rready                ,
  output             eth_axi_rvalid                ,
  output [  63:   0] eth_axi_rdata                 ,
  output [   1:   0] eth_axi_rresp                 ,
  output             eth_axi_rlast                 ,
  input              eth_axi_awvalid               ,
  output             eth_axi_awready               ,
  input  [  31:   0] eth_axi_awaddr                ,
  input  [   7:   0] eth_axi_awlen                 ,
  input  [   2:   0] eth_axi_awsize                ,
  input  [   1:   0] eth_axi_awburst               ,
  input              eth_axi_awlock                ,
  input  [   3:   0] eth_axi_awcache               ,
  input  [   2:   0] eth_axi_awprot                ,
  input              eth_axi_bready                ,
  output             eth_axi_bvalid                ,
  output [   1:   0] eth_axi_bresp                 ,
  output             eth_axi_wready                ,
  input              eth_axi_wvalid                ,
  input  [  63:   0] eth_axi_wdata                 ,
  input  [   7:   0] eth_axi_wstrb                 ,
  input              eth_axi_wlast                 ,
  output             biu2iram_icb_cmd_valid        ,
  input              biu2iram_icb_cmd_ready        ,
  output             biu2iram_icb_cmd_sel          ,
  output             biu2iram_icb_cmd_read         ,
  output [  15:   0] biu2iram_icb_cmd_addr         ,
  output [  63:   0] biu2iram_icb_cmd_wdata        ,
  output [   7:   0] biu2iram_icb_cmd_wmask        ,
  output [   2:   0] biu2iram_icb_cmd_size         ,
  output             biu2iram_icb_cmd_lock         ,
  output             biu2iram_icb_cmd_excl         ,
  output [   7:   0] biu2iram_icb_cmd_xlen         ,
  output [   1:   0] biu2iram_icb_cmd_xburst       ,
  output [   1:   0] biu2iram_icb_cmd_modes        ,
  output             biu2iram_icb_cmd_dmode        ,
  output [   2:   0] biu2iram_icb_cmd_attri        ,
  output [   1:   0] biu2iram_icb_cmd_beat         ,
  output             biu2iram_icb_rsp_ready        ,
  input              biu2iram_icb_rsp_valid        ,
  input              biu2iram_icb_rsp_err          ,
  input              biu2iram_icb_rsp_excl_ok      ,
  input  [  63:   0] biu2iram_icb_rsp_rdata        ,
  output             biu2dram_icb_cmd_valid        ,
  input              biu2dram_icb_cmd_ready        ,
  output             biu2dram_icb_cmd_sel          ,
  output             biu2dram_icb_cmd_read         ,
  output [  15:   0] biu2dram_icb_cmd_addr         ,
  output [  63:   0] biu2dram_icb_cmd_wdata        ,
  output [   7:   0] biu2dram_icb_cmd_wmask        ,
  output [   2:   0] biu2dram_icb_cmd_size         ,
  output             biu2dram_icb_cmd_lock         ,
  output             biu2dram_icb_cmd_excl         ,
  output [   7:   0] biu2dram_icb_cmd_xlen         ,
  output [   1:   0] biu2dram_icb_cmd_xburst       ,
  output [   1:   0] biu2dram_icb_cmd_modes        ,
  output             biu2dram_icb_cmd_dmode        ,
  output [   2:   0] biu2dram_icb_cmd_attri        ,
  output [   1:   0] biu2dram_icb_cmd_beat         ,
  output             biu2dram_icb_rsp_ready        ,
  input              biu2dram_icb_rsp_valid        ,
  input              biu2dram_icb_rsp_err          ,
  input              biu2dram_icb_rsp_excl_ok      ,
  input  [  63:   0] biu2dram_icb_rsp_rdata        ,
  output             addr0_icb_cmd_valid           ,
  input              addr0_icb_cmd_ready           ,
  output             addr0_icb_cmd_sel             ,
  output             addr0_icb_cmd_read            ,
  output [  31:   0] addr0_icb_cmd_addr            ,
  output [  31:   0] addr0_icb_cmd_wdata           ,
  output [   3:   0] addr0_icb_cmd_wmask           ,
  output [   2:   0] addr0_icb_cmd_size            ,
  output             addr0_icb_cmd_lock            ,
  output             addr0_icb_cmd_excl            ,
  output [   7:   0] addr0_icb_cmd_xlen            ,
  output [   1:   0] addr0_icb_cmd_xburst          ,
  output [   1:   0] addr0_icb_cmd_modes           ,
  output             addr0_icb_cmd_dmode           ,
  output [   2:   0] addr0_icb_cmd_attri           ,
  output [   1:   0] addr0_icb_cmd_beat            ,
  output             addr0_icb_rsp_ready           ,
  input              addr0_icb_rsp_valid           ,
  input              addr0_icb_rsp_err             ,
  input              addr0_icb_rsp_excl_ok         ,
  input  [  31:   0] addr0_icb_rsp_rdata           ,
  output             qspi0_ro_icb_cmd_valid        ,
  input              qspi0_ro_icb_cmd_ready        ,
  output             qspi0_ro_icb_cmd_sel          ,
  output             qspi0_ro_icb_cmd_read         ,
  output [  31:   0] qspi0_ro_icb_cmd_addr         ,
  output [  31:   0] qspi0_ro_icb_cmd_wdata        ,
  output [   3:   0] qspi0_ro_icb_cmd_wmask        ,
  output [   2:   0] qspi0_ro_icb_cmd_size         ,
  output             qspi0_ro_icb_cmd_lock         ,
  output             qspi0_ro_icb_cmd_excl         ,
  output [   7:   0] qspi0_ro_icb_cmd_xlen         ,
  output [   1:   0] qspi0_ro_icb_cmd_xburst       ,
  output [   1:   0] qspi0_ro_icb_cmd_modes        ,
  output             qspi0_ro_icb_cmd_dmode        ,
  output [   2:   0] qspi0_ro_icb_cmd_attri        ,
  output [   1:   0] qspi0_ro_icb_cmd_beat         ,
  output             qspi0_ro_icb_rsp_ready        ,
  input              qspi0_ro_icb_rsp_valid        ,
  input              qspi0_ro_icb_rsp_err          ,
  input              qspi0_ro_icb_rsp_excl_ok      ,
  input  [  31:   0] qspi0_ro_icb_rsp_rdata        ,
  output [  11:   0] eth_cfg_apb_paddr             ,
  output             eth_cfg_apb_pwrite            ,
  output             eth_cfg_apb_psel              ,
  output [   2:   0] eth_cfg_apb_pprot             ,
  output [   3:   0] eth_cfg_apb_pstrobe           ,
  output             eth_cfg_apb_penable           ,
  output [  31:   0] eth_cfg_apb_pwdata            ,
  input  [  31:   0] eth_cfg_apb_prdata            ,
  input              eth_cfg_apb_pready            ,
  input              eth_cfg_apb_pslverr           ,
  output             biu2ppi_icb_cmd_valid         ,
  input              biu2ppi_icb_cmd_ready         ,
  output             biu2ppi_icb_cmd_sel           ,
  output             biu2ppi_icb_cmd_read          ,
  output [  31:   0] biu2ppi_icb_cmd_addr          ,
  output [  31:   0] biu2ppi_icb_cmd_wdata         ,
  output [   3:   0] biu2ppi_icb_cmd_wmask         ,
  output [   2:   0] biu2ppi_icb_cmd_size          ,
  output             biu2ppi_icb_cmd_lock          ,
  output             biu2ppi_icb_cmd_excl          ,
  output [   7:   0] biu2ppi_icb_cmd_xlen          ,
  output [   1:   0] biu2ppi_icb_cmd_xburst        ,
  output [   1:   0] biu2ppi_icb_cmd_modes         ,
  output             biu2ppi_icb_cmd_dmode         ,
  output [   2:   0] biu2ppi_icb_cmd_attri         ,
  output [   1:   0] biu2ppi_icb_cmd_beat          ,
  output             biu2ppi_icb_rsp_ready         ,
  input              biu2ppi_icb_rsp_valid         ,
  input              biu2ppi_icb_rsp_err           ,
  input              biu2ppi_icb_rsp_excl_ok       ,
  input  [  31:   0] biu2ppi_icb_rsp_rdata         ,
  output             o0_axi_arvalid                ,
  input              o0_axi_arready                ,
  output [  31:   0] o0_axi_araddr                 ,
  output [   7:   0] o0_axi_arlen                  ,
  output [   2:   0] o0_axi_arsize                 ,
  output [   1:   0] o0_axi_arburst                ,
  output             o0_axi_arlock                 ,
  output [   3:   0] o0_axi_arcache                ,
  output [   2:   0] o0_axi_arprot                 ,
  output             o0_axi_rready                 ,
  input              o0_axi_rvalid                 ,
  input  [  63:   0] o0_axi_rdata                  ,
  input  [   1:   0] o0_axi_rresp                  ,
  input              o0_axi_rlast                  ,
  output             o0_axi_awvalid                ,
  input              o0_axi_awready                ,
  output [  31:   0] o0_axi_awaddr                 ,
  output [   7:   0] o0_axi_awlen                  ,
  output [   2:   0] o0_axi_awsize                 ,
  output [   1:   0] o0_axi_awburst                ,
  output             o0_axi_awlock                 ,
  output [   3:   0] o0_axi_awcache                ,
  output [   2:   0] o0_axi_awprot                 ,
  output             o0_axi_bready                 ,
  input              o0_axi_bvalid                 ,
  input  [   1:   0] o0_axi_bresp                  ,
  input              o0_axi_wready                 ,
  output             o0_axi_wvalid                 ,
  output [  63:   0] o0_axi_wdata                  ,
  output [   7:   0] o0_axi_wstrb                  ,
  output             o0_axi_wlast                  ,
  output             dummy_slv_icb_cmd_valid       ,
  input              dummy_slv_icb_cmd_ready       ,
  output             dummy_slv_icb_cmd_sel         ,
  output             dummy_slv_icb_cmd_read        ,
  output [  31:   0] dummy_slv_icb_cmd_addr        ,
  output [  63:   0] dummy_slv_icb_cmd_wdata       ,
  output [   7:   0] dummy_slv_icb_cmd_wmask       ,
  output [   2:   0] dummy_slv_icb_cmd_size        ,
  output             dummy_slv_icb_cmd_lock        ,
  output             dummy_slv_icb_cmd_excl        ,
  output [   7:   0] dummy_slv_icb_cmd_xlen        ,
  output [   1:   0] dummy_slv_icb_cmd_xburst      ,
  output [   1:   0] dummy_slv_icb_cmd_modes       ,
  output             dummy_slv_icb_cmd_dmode       ,
  output [   2:   0] dummy_slv_icb_cmd_attri       ,
  output [   1:   0] dummy_slv_icb_cmd_beat        ,
  output             dummy_slv_icb_rsp_ready       ,
  input              dummy_slv_icb_rsp_valid       ,
  input              dummy_slv_icb_rsp_err         ,
  input              dummy_slv_icb_rsp_excl_ok     ,
  input  [  63:   0] dummy_slv_icb_rsp_rdata       ,
  input  [   2:   0] i_axi_aruser                  ,
  output [   2:   0] i_axi_ruser                   ,
  input  [   2:   0] i_axi_arid                    ,
  output [   2:   0] i_axi_rid                     ,
  input  [   2:   0] i_axi_awuser                  ,
  output [   2:   0] i_axi_buser                   ,
  input  [   2:   0] i_axi_awid                    ,
  output [   2:   0] i_axi_bid                     ,
  input  [   2:   0] dummy_axi_arid                ,
  output [   2:   0] dummy_axi_rid                 ,
  input  [   2:   0] dummy_axi_awid                ,
  output [   2:   0] dummy_axi_bid                 ,
  input              eth_axi_clk                   ,
  input              eth_axi_rst_n                 ,
  input              biu2iram_icb_clk_en           ,
  input              biu2iram_icb_clk              ,
  input              biu2iram_icb_rst_n            ,
  input              biu2dram_icb_clk_en           ,
  input              biu2dram_icb_clk              ,
  input              biu2dram_icb_rst_n            ,
  input              o0_axi_clk                    ,
  input              o0_axi_rst_n                  ,
  output [   2:   0] o0_axi_arid                   ,
  input  [   2:   0] o0_axi_rid                    ,
  output [   2:   0] o0_axi_awid                   ,
  input  [   2:   0] o0_axi_bid                    ,
  input              clkgate_bypass                ,
  input              clk                           ,
  input              rst_n                         
  );
  wire clk_fab;
  localparam PAYLOAD_NORST = 0 ;
  localparam RSP_CHECK_CMD_OUTS  = 1;
  localparam RRBIN_CUT_TIMING = 1;
  localparam CLKGATE_PARAM = 1;
  localparam SUPPORT_W2N_ID_OOO = 0;
  wire fab_active;
  generate
  if(CLKGATE_PARAM == 1) begin: clkgate_gen
      e603_clkgate u_fab_clkgate(
        .clk_in   (clk),
        .clkgate_bypass(clkgate_bypass  ),
        .clock_en (fab_active),
        .clk_out  (clk_fab)
      );
  end
  else begin: no_clkgate_gen
    assign clk_fab = clk;
  end
  endgenerate
               wire eth_axi_rst_n_sync_4port;
               wire eth_axi_rst_n_sync_4fab;
               wire eth_axi_rst_n_sync_i = eth_axi_rst_n & rst_n;
  e603_reset_sync u_eth_axi__rst_sync_4port(
    .clk      (eth_axi_clk), 
    .rst_n_a  (eth_axi_rst_n_sync_i),
    .reset_bypass(clkgate_bypass), 
    .rst_n_sync(eth_axi_rst_n_sync_4port)
  );
  e603_reset_sync u_eth_axi__rst_sync_4fab(
    .clk      (clk), 
    .rst_n_a  (eth_axi_rst_n_sync_i),
    .reset_bypass(clkgate_bypass), 
    .rst_n_sync(eth_axi_rst_n_sync_4fab)
  );
               wire o0_axi_rst_n_sync_4port;
               wire o0_axi_rst_n_sync_4fab;
               wire o0_axi_rst_n_sync_i = o0_axi_rst_n & rst_n;
  e603_reset_sync u_o0_axi__rst_sync_4port(
    .clk      (o0_axi_clk), 
    .rst_n_a  (o0_axi_rst_n_sync_i),
    .reset_bypass(clkgate_bypass), 
    .rst_n_sync(o0_axi_rst_n_sync_4port)
  );
  e603_reset_sync u_o0_axi__rst_sync_4fab(
    .clk      (clk), 
    .rst_n_a  (o0_axi_rst_n_sync_i),
    .reset_bypass(clkgate_bypass), 
    .rst_n_sync(o0_axi_rst_n_sync_4fab)
  );
      wire                mst_grp_0_ro_icb_cmd_valid    ;
  wire                mst_grp_0_ro_icb_cmd_ready    ;
  wire                mst_grp_0_ro_icb_cmd_sel      ;
  wire                mst_grp_0_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_0_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_0_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_0_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_0_ro_icb_cmd_size     ;
  wire                mst_grp_0_ro_icb_cmd_lock     ;
  wire                mst_grp_0_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_0_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_0_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_0_ro_icb_cmd_modes    ;
  wire                mst_grp_0_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_0_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_0_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_0_ro_icb_cmd_usr      ;
  wire                mst_grp_0_ro_icb_rsp_ready    ;
  wire                mst_grp_0_ro_icb_rsp_valid    ;
  wire                mst_grp_0_ro_icb_rsp_err      ;
  wire                mst_grp_0_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_0_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_0_ro_icb_rsp_usr      ;
      wire                mst_grp_0_wo_icb_cmd_valid    ;
  wire                mst_grp_0_wo_icb_cmd_ready    ;
  wire                mst_grp_0_wo_icb_cmd_sel      ;
  wire                mst_grp_0_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_0_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_0_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_0_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_0_wo_icb_cmd_size     ;
  wire                mst_grp_0_wo_icb_cmd_lock     ;
  wire                mst_grp_0_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_0_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_0_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_0_wo_icb_cmd_modes    ;
  wire                mst_grp_0_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_0_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_0_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_0_wo_icb_cmd_usr      ;
  wire                mst_grp_0_wo_icb_rsp_ready    ;
  wire                mst_grp_0_wo_icb_rsp_valid    ;
  wire                mst_grp_0_wo_icb_rsp_err      ;
  wire                mst_grp_0_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_0_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_0_wo_icb_rsp_usr      ;
                 wire                mst_g0_p0_icb_cmd_valid       ;
  wire                mst_g0_p0_icb_cmd_ready       ;
  wire                mst_g0_p0_icb_cmd_sel         ;
  wire                mst_g0_p0_icb_cmd_read        ;
  wire    [  31:   0] mst_g0_p0_icb_cmd_addr        ;
  wire    [  63:   0] mst_g0_p0_icb_cmd_wdata       ;
  wire    [   7:   0] mst_g0_p0_icb_cmd_wmask       ;
  wire    [   2:   0] mst_g0_p0_icb_cmd_size        ;
  wire                mst_g0_p0_icb_cmd_lock        ;
  wire                mst_g0_p0_icb_cmd_excl        ;
  wire    [   7:   0] mst_g0_p0_icb_cmd_xlen        ;
  wire    [   1:   0] mst_g0_p0_icb_cmd_xburst      ;
  wire    [   1:   0] mst_g0_p0_icb_cmd_modes       ;
  wire                mst_g0_p0_icb_cmd_dmode       ;
  wire    [   2:   0] mst_g0_p0_icb_cmd_attri       ;
  wire    [   1:   0] mst_g0_p0_icb_cmd_beat        ;
  wire    [   2:   0] mst_g0_p0_icb_cmd_usr         ;
  wire                mst_g0_p0_icb_rsp_ready       ;
  wire                mst_g0_p0_icb_rsp_valid       ;
  wire                mst_g0_p0_icb_rsp_err         ;
  wire                mst_g0_p0_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_g0_p0_icb_rsp_rdata       ;
  wire    [   2:   0] mst_g0_p0_icb_rsp_usr         ;
                wire [3-1:0] mst_g0_p0_icb_cmd_id;
                wire [3-1:0] mst_g0_p0_icb_rsp_id;
                wire                  mst_g0_p0_icb_rsp_last;
                 wire                mst_g0_p0_w2n_ro_icb_cmd_valid ;
  wire                mst_g0_p0_w2n_ro_icb_cmd_ready ;
  wire                mst_g0_p0_w2n_ro_icb_cmd_sel  ;
  wire                mst_g0_p0_w2n_ro_icb_cmd_read ;
  wire    [  31:   0] mst_g0_p0_w2n_ro_icb_cmd_addr ;
  wire    [  63:   0] mst_g0_p0_w2n_ro_icb_cmd_wdata ;
  wire    [   7:   0] mst_g0_p0_w2n_ro_icb_cmd_wmask ;
  wire    [   2:   0] mst_g0_p0_w2n_ro_icb_cmd_size ;
  wire                mst_g0_p0_w2n_ro_icb_cmd_lock ;
  wire                mst_g0_p0_w2n_ro_icb_cmd_excl ;
  wire    [   7:   0] mst_g0_p0_w2n_ro_icb_cmd_xlen ;
  wire    [   1:   0] mst_g0_p0_w2n_ro_icb_cmd_xburst ;
  wire    [   1:   0] mst_g0_p0_w2n_ro_icb_cmd_modes ;
  wire                mst_g0_p0_w2n_ro_icb_cmd_dmode ;
  wire    [   2:   0] mst_g0_p0_w2n_ro_icb_cmd_attri ;
  wire    [   1:   0] mst_g0_p0_w2n_ro_icb_cmd_beat ;
  wire    [   2:   0] mst_g0_p0_w2n_ro_icb_cmd_usr  ;
  wire                mst_g0_p0_w2n_ro_icb_rsp_ready ;
  wire                mst_g0_p0_w2n_ro_icb_rsp_valid ;
  wire                mst_g0_p0_w2n_ro_icb_rsp_err  ;
  wire                mst_g0_p0_w2n_ro_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g0_p0_w2n_ro_icb_rsp_rdata ;
  wire    [   2:   0] mst_g0_p0_w2n_ro_icb_rsp_usr  ;
                 wire                mst_g0_p0_w2n_wo_icb_cmd_valid ;
  wire                mst_g0_p0_w2n_wo_icb_cmd_ready ;
  wire                mst_g0_p0_w2n_wo_icb_cmd_sel  ;
  wire                mst_g0_p0_w2n_wo_icb_cmd_read ;
  wire    [  31:   0] mst_g0_p0_w2n_wo_icb_cmd_addr ;
  wire    [  63:   0] mst_g0_p0_w2n_wo_icb_cmd_wdata ;
  wire    [   7:   0] mst_g0_p0_w2n_wo_icb_cmd_wmask ;
  wire    [   2:   0] mst_g0_p0_w2n_wo_icb_cmd_size ;
  wire                mst_g0_p0_w2n_wo_icb_cmd_lock ;
  wire                mst_g0_p0_w2n_wo_icb_cmd_excl ;
  wire    [   7:   0] mst_g0_p0_w2n_wo_icb_cmd_xlen ;
  wire    [   1:   0] mst_g0_p0_w2n_wo_icb_cmd_xburst ;
  wire    [   1:   0] mst_g0_p0_w2n_wo_icb_cmd_modes ;
  wire                mst_g0_p0_w2n_wo_icb_cmd_dmode ;
  wire    [   2:   0] mst_g0_p0_w2n_wo_icb_cmd_attri ;
  wire    [   1:   0] mst_g0_p0_w2n_wo_icb_cmd_beat ;
  wire    [   2:   0] mst_g0_p0_w2n_wo_icb_cmd_usr  ;
  wire                mst_g0_p0_w2n_wo_icb_rsp_ready ;
  wire                mst_g0_p0_w2n_wo_icb_rsp_valid ;
  wire                mst_g0_p0_w2n_wo_icb_rsp_err  ;
  wire                mst_g0_p0_w2n_wo_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g0_p0_w2n_wo_icb_rsp_rdata ;
  wire    [   2:   0] mst_g0_p0_w2n_wo_icb_rsp_usr  ;
    wire i_axi_bus_active;
                 wire                mst_g0_p0_ro_icb_cmd_valid    ;
  wire                mst_g0_p0_ro_icb_cmd_ready    ;
  wire                mst_g0_p0_ro_icb_cmd_sel      ;
  wire                mst_g0_p0_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_g0_p0_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_g0_p0_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_g0_p0_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_g0_p0_ro_icb_cmd_size     ;
  wire                mst_g0_p0_ro_icb_cmd_lock     ;
  wire                mst_g0_p0_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_g0_p0_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_g0_p0_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_g0_p0_ro_icb_cmd_modes    ;
  wire                mst_g0_p0_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_g0_p0_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_g0_p0_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_g0_p0_ro_icb_cmd_usr      ;
  wire                mst_g0_p0_ro_icb_rsp_ready    ;
  wire                mst_g0_p0_ro_icb_rsp_valid    ;
  wire                mst_g0_p0_ro_icb_rsp_err      ;
  wire                mst_g0_p0_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_g0_p0_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_g0_p0_ro_icb_rsp_usr      ;
                    wire [3-1:0] mst_g0_p0_ro_icb_cmd_id;
                    wire [3-1:0] mst_g0_p0_ro_icb_rsp_id;
                    wire                  mst_g0_p0_ro_icb_rsp_last;
    wire mst_g0_p0_ro_icb_bus_active;
                              wire[3-1:0] mst_g0_p0_ro_icb_cmd_usr_pre;
               assign mst_g0_p0_ro_icb_cmd_usr = mst_g0_p0_ro_icb_cmd_usr_pre;
  e603_subsys_gnrl_axi2ficb_read_id # (
      .ALLOW_FIX_BURST(1),
      .ID_W(3),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .RATIO_FIFO_DP(2),
      .AW(32),
      .DW(64), 
      .MW(64/8), 
      .FIFO_OUTS_NUM (128),
      .USR_W (3)
    )u_i_axi_axi2ficb_read(
  .reset_flag_r  (1'b0),
  .axi_bus_clk_en(1'b1),
  .icb_clk_en(1'b1),
      .axi_arvalid                    (i_axi_arvalid                            ),
  .axi_arready                    (i_axi_arready                            ),
  .axi_arlen                      (i_axi_arlen                   [   7:   0]),
  .axi_arsize                     (i_axi_arsize                  [   2:   0]),
  .axi_arburst                    (i_axi_arburst                 [   1:   0]),
  .axi_arlock                     (i_axi_arlock                             ),
  .axi_arcache                    (i_axi_arcache                 [   3:   0]),
  .axi_arprot                     (i_axi_arprot                  [   2:   0]),
  .axi_rready                     (i_axi_rready                             ),
  .axi_rvalid                     (i_axi_rvalid                             ),
  .axi_rdata                      (i_axi_rdata                   [  63:   0]),
  .axi_rresp                      (i_axi_rresp                   [   1:   0]),
  .axi_rlast                      (i_axi_rlast                              ),
      .axi_araddr(i_axi_araddr[32-1:0]),
      .axi_aruser(i_axi_aruser),
      .axi_ruser(i_axi_ruser),
      .axi_arid(i_axi_arid),
      .axi_rid (i_axi_rid ),
        .icb_rcmd_valid                 (mst_g0_p0_ro_icb_cmd_valid               ),
  .icb_rcmd_ready                 (mst_g0_p0_ro_icb_cmd_ready               ),
  .icb_rcmd_sel                   (mst_g0_p0_ro_icb_cmd_sel                 ),
  .icb_rcmd_read                  (mst_g0_p0_ro_icb_cmd_read                ),
  .icb_rcmd_addr                  (mst_g0_p0_ro_icb_cmd_addr     [  31:   0]),
  .icb_rcmd_wdata                 (mst_g0_p0_ro_icb_cmd_wdata    [  63:   0]),
  .icb_rcmd_wmask                 (mst_g0_p0_ro_icb_cmd_wmask    [   7:   0]),
  .icb_rcmd_size                  (mst_g0_p0_ro_icb_cmd_size     [   2:   0]),
  .icb_rcmd_excl                  (mst_g0_p0_ro_icb_cmd_excl                ),
  .icb_rcmd_xlen                  (mst_g0_p0_ro_icb_cmd_xlen     [   7:   0]),
  .icb_rcmd_xburst                (mst_g0_p0_ro_icb_cmd_xburst   [   1:   0]),
  .icb_rcmd_modes                 (mst_g0_p0_ro_icb_cmd_modes    [   1:   0]),
  .icb_rcmd_dmode                 (mst_g0_p0_ro_icb_cmd_dmode               ),
  .icb_rcmd_attri                 (mst_g0_p0_ro_icb_cmd_attri    [   2:   0]),
  .icb_rcmd_beat                  (mst_g0_p0_ro_icb_cmd_beat     [   1:   0]),
  .icb_rrsp_ready                 (mst_g0_p0_ro_icb_rsp_ready               ),
  .icb_rrsp_valid                 (mst_g0_p0_ro_icb_rsp_valid               ),
  .icb_rrsp_err                   (mst_g0_p0_ro_icb_rsp_err                 ),
  .icb_rrsp_excl_ok               (mst_g0_p0_ro_icb_rsp_excl_ok             ),
  .icb_rrsp_rdata                 (mst_g0_p0_ro_icb_rsp_rdata    [  63:   0]),
      .icb_rcmd_usr(mst_g0_p0_ro_icb_cmd_usr_pre),
      .icb_rrsp_usr(mst_g0_p0_ro_icb_rsp_usr[3-1:0]),
      .icb_rcmd_id(mst_g0_p0_ro_icb_cmd_id),
      .icb_rrsp_id(mst_g0_p0_ro_icb_rsp_id),
      .icb_rrsp_last(mst_g0_p0_ro_icb_rsp_last),
      .axi2icb_read_active (mst_g0_p0_ro_icb_bus_active),
      .clk  (clk_fab),  
      .rst_n(rst_n)
    );
    assign mst_g0_p0_ro_icb_cmd_lock = 1'b0;
                 wire                mst_g0_p0_wo_icb_cmd_valid    ;
  wire                mst_g0_p0_wo_icb_cmd_ready    ;
  wire                mst_g0_p0_wo_icb_cmd_sel      ;
  wire                mst_g0_p0_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_g0_p0_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_g0_p0_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_g0_p0_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_g0_p0_wo_icb_cmd_size     ;
  wire                mst_g0_p0_wo_icb_cmd_lock     ;
  wire                mst_g0_p0_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_g0_p0_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_g0_p0_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_g0_p0_wo_icb_cmd_modes    ;
  wire                mst_g0_p0_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_g0_p0_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_g0_p0_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_g0_p0_wo_icb_cmd_usr      ;
  wire                mst_g0_p0_wo_icb_rsp_ready    ;
  wire                mst_g0_p0_wo_icb_rsp_valid    ;
  wire                mst_g0_p0_wo_icb_rsp_err      ;
  wire                mst_g0_p0_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_g0_p0_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_g0_p0_wo_icb_rsp_usr      ;
                    wire [3-1:0] mst_g0_p0_wo_icb_cmd_id;
                    wire [3-1:0] mst_g0_p0_wo_icb_rsp_id;
                    wire                  mst_g0_p0_wo_icb_rsp_last;
    wire mst_g0_p0_wo_icb_bus_active;
                              wire[3-1:0] mst_g0_p0_wo_icb_cmd_usr_pre;
               assign mst_g0_p0_wo_icb_cmd_usr = mst_g0_p0_wo_icb_cmd_usr_pre;
  e603_subsys_gnrl_axi2ficb_write_id # (
      .ALLOW_FIX_BURST(1),
      .ID_W(3),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .RATIO_FIFO_DP(2),
      .AW(32),
      .DW(64), 
      .MW(64/8), 
      .FIFO_OUTS_NUM (128),
      .USR_W (3)
    )u_mst_g0_p0_wo_icb_axi2ficb_write(
  .reset_flag_r  (1'b0),
  .axi_bus_clk_en(1'b1),
  .icb_clk_en(1'b1),
      .axi_awvalid                    (i_axi_awvalid                            ),
  .axi_awready                    (i_axi_awready                            ),
  .axi_awlen                      (i_axi_awlen                   [   7:   0]),
  .axi_awsize                     (i_axi_awsize                  [   2:   0]),
  .axi_awburst                    (i_axi_awburst                 [   1:   0]),
  .axi_awlock                     (i_axi_awlock                             ),
  .axi_awcache                    (i_axi_awcache                 [   3:   0]),
  .axi_awprot                     (i_axi_awprot                  [   2:   0]),
  .axi_bready                     (i_axi_bready                             ),
  .axi_bvalid                     (i_axi_bvalid                             ),
  .axi_bresp                      (i_axi_bresp                   [   1:   0]),
  .axi_wready                     (i_axi_wready                             ),
  .axi_wvalid                     (i_axi_wvalid                             ),
  .axi_wdata                      (i_axi_wdata                   [  63:   0]),
  .axi_wstrb                      (i_axi_wstrb                   [   7:   0]),
  .axi_wlast                      (i_axi_wlast                              ),
      .axi_awaddr(i_axi_awaddr[32-1:0]),
      .axi_awuser(i_axi_awuser),
      .axi_buser(i_axi_buser),
      .axi_awid(i_axi_awid),
      .axi_bid (i_axi_bid ),
        .icb_wcmd_valid                 (mst_g0_p0_wo_icb_cmd_valid               ),
  .icb_wcmd_ready                 (mst_g0_p0_wo_icb_cmd_ready               ),
  .icb_wcmd_sel                   (mst_g0_p0_wo_icb_cmd_sel                 ),
  .icb_wcmd_read                  (mst_g0_p0_wo_icb_cmd_read                ),
  .icb_wcmd_addr                  (mst_g0_p0_wo_icb_cmd_addr     [  31:   0]),
  .icb_wcmd_wdata                 (mst_g0_p0_wo_icb_cmd_wdata    [  63:   0]),
  .icb_wcmd_wmask                 (mst_g0_p0_wo_icb_cmd_wmask    [   7:   0]),
  .icb_wcmd_size                  (mst_g0_p0_wo_icb_cmd_size     [   2:   0]),
  .icb_wcmd_lock                  (mst_g0_p0_wo_icb_cmd_lock                ),
  .icb_wcmd_excl                  (mst_g0_p0_wo_icb_cmd_excl                ),
  .icb_wcmd_xlen                  (mst_g0_p0_wo_icb_cmd_xlen     [   7:   0]),
  .icb_wcmd_xburst                (mst_g0_p0_wo_icb_cmd_xburst   [   1:   0]),
  .icb_wcmd_modes                 (mst_g0_p0_wo_icb_cmd_modes    [   1:   0]),
  .icb_wcmd_dmode                 (mst_g0_p0_wo_icb_cmd_dmode               ),
  .icb_wcmd_attri                 (mst_g0_p0_wo_icb_cmd_attri    [   2:   0]),
  .icb_wcmd_beat                  (mst_g0_p0_wo_icb_cmd_beat     [   1:   0]),
  .icb_wrsp_ready                 (mst_g0_p0_wo_icb_rsp_ready               ),
  .icb_wrsp_valid                 (mst_g0_p0_wo_icb_rsp_valid               ),
  .icb_wrsp_err                   (mst_g0_p0_wo_icb_rsp_err                 ),
  .icb_wrsp_excl_ok               (mst_g0_p0_wo_icb_rsp_excl_ok             ),
      .icb_wcmd_usr(mst_g0_p0_wo_icb_cmd_usr_pre),
      .icb_wrsp_usr(mst_g0_p0_wo_icb_rsp_usr[3-1:0]),
      .icb_wcmd_id(mst_g0_p0_wo_icb_cmd_id),
      .icb_wrsp_id(mst_g0_p0_wo_icb_rsp_id),
      .axi2icb_write_active (mst_g0_p0_wo_icb_bus_active),
      .clk  (clk_fab),  
      .rst_n(rst_n)
    );
   assign i_axi_bus_active = 1'b0
                     | mst_g0_p0_ro_icb_bus_active
                     | mst_g0_p0_wo_icb_bus_active
                 ;
   wire mst_g0_p0_ro_icb_id_gen_ready;
   wire [1:0] mst_g0_p0_ro_icb_cmd_beat_raw;
   wire [7:0] mst_g0_p0_ro_icb_cmd_xlen_raw;
   e603_subsys_gnrl_ficb_id_gen # (
     .OUTS_FIFO_DP (128+1),
     .ID_W         (3)
   ) u_mst_g0_p0_ro_icb_ficb_id_gen(
     .i_icb_cmd_valid(mst_g0_p0_ro_icb_cmd_valid), 
     .i_icb_cmd_ready(mst_g0_p0_ro_icb_cmd_ready), 
     .i_icb_cmd_id   (mst_g0_p0_ro_icb_cmd_id),
     .i_icb_cmd_xburst (mst_g0_p0_ro_icb_cmd_xburst),
     .i_icb_cmd_beat   (mst_g0_p0_ro_icb_cmd_beat),
     .i_icb_cmd_xlen   (mst_g0_p0_ro_icb_cmd_xlen),
     .i_icb_cmd_size   (mst_g0_p0_ro_icb_cmd_size),
     .o_icb_cmd_beat   (mst_g0_p0_ro_icb_cmd_beat_raw),
     .o_icb_cmd_xlen   (mst_g0_p0_ro_icb_cmd_xlen_raw),
     .ficb_id_gen_ready (mst_g0_p0_ro_icb_id_gen_ready),
     .i_icb_rsp_valid(mst_g0_p0_ro_icb_rsp_valid), 
     .i_icb_rsp_ready(mst_g0_p0_ro_icb_rsp_ready), 
     .i_icb_rsp_id   (mst_g0_p0_ro_icb_rsp_id),
     .i_icb_rsp_last   (mst_g0_p0_ro_icb_rsp_last),
    .clk  (clk_fab),  
    .rst_n(rst_n)
     );
    wire mst_g0_p0_ro_icb_cmd_valid_raw;
    wire mst_g0_p0_ro_icb_cmd_ready_raw;
    assign mst_g0_p0_ro_icb_cmd_valid_raw = (mst_g0_p0_ro_icb_id_gen_ready) & mst_g0_p0_ro_icb_cmd_valid;
    assign mst_g0_p0_ro_icb_cmd_ready     = (mst_g0_p0_ro_icb_id_gen_ready) & mst_g0_p0_ro_icb_cmd_ready_raw;
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (128),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g0_p0_ro_icb_ficb_wconv(
      .i_icb_cmd_read(1'b1),
                .i_icb_cmd_wdata (64'b0),
                .i_icb_cmd_wmask (8'b0),
                .i_icb_cmd_valid(mst_g0_p0_ro_icb_cmd_valid_raw),
                .i_icb_cmd_ready(mst_g0_p0_ro_icb_cmd_ready_raw),
                .i_icb_cmd_beat (mst_g0_p0_ro_icb_cmd_beat_raw),
                .i_icb_cmd_xlen (mst_g0_p0_ro_icb_cmd_xlen_raw),
        .i_icb_cmd_sel                  (mst_g0_p0_ro_icb_cmd_sel                 ),
  .i_icb_cmd_addr                 (mst_g0_p0_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_size                 (mst_g0_p0_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_g0_p0_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_g0_p0_ro_icb_cmd_excl                ),
  .i_icb_cmd_xburst               (mst_g0_p0_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_g0_p0_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_g0_p0_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_g0_p0_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_usr                  (mst_g0_p0_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_g0_p0_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_g0_p0_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_g0_p0_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_g0_p0_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_g0_p0_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_g0_p0_ro_icb_rsp_usr      [   2:   0]),
        .o_icb_cmd_valid                (mst_g0_p0_w2n_ro_icb_cmd_valid            ),
  .o_icb_cmd_ready                (mst_g0_p0_w2n_ro_icb_cmd_ready            ),
  .o_icb_cmd_sel                  (mst_g0_p0_w2n_ro_icb_cmd_sel             ),
  .o_icb_cmd_read                 (mst_g0_p0_w2n_ro_icb_cmd_read            ),
  .o_icb_cmd_addr                 (mst_g0_p0_w2n_ro_icb_cmd_addr [  31:   0]),
  .o_icb_cmd_wdata                (mst_g0_p0_w2n_ro_icb_cmd_wdata [  63:   0]),
  .o_icb_cmd_wmask                (mst_g0_p0_w2n_ro_icb_cmd_wmask [   7:   0]),
  .o_icb_cmd_size                 (mst_g0_p0_w2n_ro_icb_cmd_size [   2:   0]),
  .o_icb_cmd_lock                 (mst_g0_p0_w2n_ro_icb_cmd_lock            ),
  .o_icb_cmd_excl                 (mst_g0_p0_w2n_ro_icb_cmd_excl            ),
  .o_icb_cmd_xlen                 (mst_g0_p0_w2n_ro_icb_cmd_xlen [   7:   0]),
  .o_icb_cmd_xburst               (mst_g0_p0_w2n_ro_icb_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (mst_g0_p0_w2n_ro_icb_cmd_modes [   1:   0]),
  .o_icb_cmd_dmode                (mst_g0_p0_w2n_ro_icb_cmd_dmode            ),
  .o_icb_cmd_attri                (mst_g0_p0_w2n_ro_icb_cmd_attri [   2:   0]),
  .o_icb_cmd_beat                 (mst_g0_p0_w2n_ro_icb_cmd_beat [   1:   0]),
  .o_icb_cmd_usr                  (mst_g0_p0_w2n_ro_icb_cmd_usr  [   2:   0]),
  .o_icb_rsp_ready                (mst_g0_p0_w2n_ro_icb_rsp_ready            ),
  .o_icb_rsp_valid                (mst_g0_p0_w2n_ro_icb_rsp_valid            ),
  .o_icb_rsp_err                  (mst_g0_p0_w2n_ro_icb_rsp_err             ),
  .o_icb_rsp_excl_ok              (mst_g0_p0_w2n_ro_icb_rsp_excl_ok            ),
  .o_icb_rsp_rdata                (mst_g0_p0_w2n_ro_icb_rsp_rdata [  63:   0]),
  .o_icb_rsp_usr                  (mst_g0_p0_w2n_ro_icb_rsp_usr  [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   wire mst_g0_p0_wo_icb_id_gen_ready;
   wire [1:0] mst_g0_p0_wo_icb_cmd_beat_raw;
   wire [7:0] mst_g0_p0_wo_icb_cmd_xlen_raw;
   e603_subsys_gnrl_ficb_id_gen # (
     .OUTS_FIFO_DP (128+1),
     .ID_W         (3)
   ) u_mst_g0_p0_wo_icb_ficb_id_gen(
     .i_icb_cmd_valid(mst_g0_p0_wo_icb_cmd_valid), 
     .i_icb_cmd_ready(mst_g0_p0_wo_icb_cmd_ready), 
     .i_icb_cmd_id   (mst_g0_p0_wo_icb_cmd_id),
     .i_icb_cmd_xburst (mst_g0_p0_wo_icb_cmd_xburst),
     .i_icb_cmd_beat   (mst_g0_p0_wo_icb_cmd_beat),
     .i_icb_cmd_xlen   (mst_g0_p0_wo_icb_cmd_xlen),
     .i_icb_cmd_size   (mst_g0_p0_wo_icb_cmd_size),
     .o_icb_cmd_beat   (mst_g0_p0_wo_icb_cmd_beat_raw),
     .o_icb_cmd_xlen   (mst_g0_p0_wo_icb_cmd_xlen_raw),
     .ficb_id_gen_ready (mst_g0_p0_wo_icb_id_gen_ready),
     .i_icb_rsp_valid(mst_g0_p0_wo_icb_rsp_valid), 
     .i_icb_rsp_ready(mst_g0_p0_wo_icb_rsp_ready), 
     .i_icb_rsp_id   (mst_g0_p0_wo_icb_rsp_id),
     .i_icb_rsp_last   (mst_g0_p0_wo_icb_rsp_last),
    .clk  (clk_fab),  
    .rst_n(rst_n)
     );
    wire mst_g0_p0_wo_icb_cmd_valid_raw;
    wire mst_g0_p0_wo_icb_cmd_ready_raw;
    assign mst_g0_p0_wo_icb_cmd_valid_raw = (mst_g0_p0_wo_icb_id_gen_ready) & mst_g0_p0_wo_icb_cmd_valid;
    assign mst_g0_p0_wo_icb_cmd_ready     = (mst_g0_p0_wo_icb_id_gen_ready) & mst_g0_p0_wo_icb_cmd_ready_raw;
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (128),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g0_p0_wo_icb_ficb_wconv(
                .i_icb_cmd_valid(mst_g0_p0_wo_icb_cmd_valid_raw),
                .i_icb_cmd_ready(mst_g0_p0_wo_icb_cmd_ready_raw),
                .i_icb_cmd_xlen (mst_g0_p0_wo_icb_cmd_xlen_raw),
                .i_icb_cmd_beat (mst_g0_p0_wo_icb_cmd_beat_raw),
        .i_icb_cmd_sel                  (mst_g0_p0_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_g0_p0_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_g0_p0_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_g0_p0_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_g0_p0_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_g0_p0_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_g0_p0_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_g0_p0_wo_icb_cmd_excl                ),
  .i_icb_cmd_xburst               (mst_g0_p0_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_g0_p0_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_g0_p0_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_g0_p0_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_usr                  (mst_g0_p0_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_g0_p0_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_g0_p0_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_g0_p0_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_g0_p0_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_g0_p0_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_g0_p0_wo_icb_rsp_usr      [   2:   0]),
                .o_icb_rsp_rdata (64'b0),
        .o_icb_cmd_valid                (mst_g0_p0_w2n_wo_icb_cmd_valid            ),
  .o_icb_cmd_ready                (mst_g0_p0_w2n_wo_icb_cmd_ready            ),
  .o_icb_cmd_sel                  (mst_g0_p0_w2n_wo_icb_cmd_sel             ),
  .o_icb_cmd_read                 (mst_g0_p0_w2n_wo_icb_cmd_read            ),
  .o_icb_cmd_addr                 (mst_g0_p0_w2n_wo_icb_cmd_addr [  31:   0]),
  .o_icb_cmd_wdata                (mst_g0_p0_w2n_wo_icb_cmd_wdata [  63:   0]),
  .o_icb_cmd_wmask                (mst_g0_p0_w2n_wo_icb_cmd_wmask [   7:   0]),
  .o_icb_cmd_size                 (mst_g0_p0_w2n_wo_icb_cmd_size [   2:   0]),
  .o_icb_cmd_lock                 (mst_g0_p0_w2n_wo_icb_cmd_lock            ),
  .o_icb_cmd_excl                 (mst_g0_p0_w2n_wo_icb_cmd_excl            ),
  .o_icb_cmd_xlen                 (mst_g0_p0_w2n_wo_icb_cmd_xlen [   7:   0]),
  .o_icb_cmd_xburst               (mst_g0_p0_w2n_wo_icb_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (mst_g0_p0_w2n_wo_icb_cmd_modes [   1:   0]),
  .o_icb_cmd_dmode                (mst_g0_p0_w2n_wo_icb_cmd_dmode            ),
  .o_icb_cmd_attri                (mst_g0_p0_w2n_wo_icb_cmd_attri [   2:   0]),
  .o_icb_cmd_beat                 (mst_g0_p0_w2n_wo_icb_cmd_beat [   1:   0]),
  .o_icb_cmd_usr                  (mst_g0_p0_w2n_wo_icb_cmd_usr  [   2:   0]),
  .o_icb_rsp_ready                (mst_g0_p0_w2n_wo_icb_rsp_ready            ),
  .o_icb_rsp_valid                (mst_g0_p0_w2n_wo_icb_rsp_valid            ),
  .o_icb_rsp_err                  (mst_g0_p0_w2n_wo_icb_rsp_err             ),
  .o_icb_rsp_excl_ok              (mst_g0_p0_w2n_wo_icb_rsp_excl_ok            ),
  .o_icb_rsp_usr                  (mst_g0_p0_w2n_wo_icb_rsp_usr  [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   e603_subsys_mgrp0_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0),
      .ICB_FIFO_RSP_DP        (0),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (128  ),
      .ARBT_FIFO_OUTS_CNT_W(8),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o0_ro_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g0_p0_w2n_ro_icb_cmd_valid            ),
  .i0_icb_cmd_ready               (mst_g0_p0_w2n_ro_icb_cmd_ready            ),
  .i0_icb_cmd_sel                 (mst_g0_p0_w2n_ro_icb_cmd_sel             ),
  .i0_icb_cmd_read                (mst_g0_p0_w2n_ro_icb_cmd_read            ),
  .i0_icb_cmd_addr                (mst_g0_p0_w2n_ro_icb_cmd_addr [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g0_p0_w2n_ro_icb_cmd_wdata [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g0_p0_w2n_ro_icb_cmd_wmask [   7:   0]),
  .i0_icb_cmd_size                (mst_g0_p0_w2n_ro_icb_cmd_size [   2:   0]),
  .i0_icb_cmd_lock                (mst_g0_p0_w2n_ro_icb_cmd_lock            ),
  .i0_icb_cmd_excl                (mst_g0_p0_w2n_ro_icb_cmd_excl            ),
  .i0_icb_cmd_xlen                (mst_g0_p0_w2n_ro_icb_cmd_xlen [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g0_p0_w2n_ro_icb_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (mst_g0_p0_w2n_ro_icb_cmd_modes [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g0_p0_w2n_ro_icb_cmd_dmode            ),
  .i0_icb_cmd_attri               (mst_g0_p0_w2n_ro_icb_cmd_attri [   2:   0]),
  .i0_icb_cmd_beat                (mst_g0_p0_w2n_ro_icb_cmd_beat [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g0_p0_w2n_ro_icb_cmd_usr  [   2:   0]),
  .i0_icb_rsp_ready               (mst_g0_p0_w2n_ro_icb_rsp_ready            ),
  .i0_icb_rsp_valid               (mst_g0_p0_w2n_ro_icb_rsp_valid            ),
  .i0_icb_rsp_err                 (mst_g0_p0_w2n_ro_icb_rsp_err             ),
  .i0_icb_rsp_excl_ok             (mst_g0_p0_w2n_ro_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g0_p0_w2n_ro_icb_rsp_rdata [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g0_p0_w2n_ro_icb_rsp_usr  [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_0_ro_icb_cmd_valid               ),
  .o_icb_cmd_ready                (mst_grp_0_ro_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (mst_grp_0_ro_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (mst_grp_0_ro_icb_cmd_read                ),
  .o_icb_cmd_addr                 (mst_grp_0_ro_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_0_ro_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_0_ro_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_0_ro_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_0_ro_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (mst_grp_0_ro_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (mst_grp_0_ro_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_0_ro_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_0_ro_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_0_ro_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (mst_grp_0_ro_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_0_ro_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_0_ro_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_0_ro_icb_rsp_ready               ),
  .o_icb_rsp_valid                (mst_grp_0_ro_icb_rsp_valid               ),
  .o_icb_rsp_err                  (mst_grp_0_ro_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (mst_grp_0_ro_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (mst_grp_0_ro_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_0_ro_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_mgrp0_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0),
      .ICB_FIFO_RSP_DP        (0),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (128  ),
      .ARBT_FIFO_OUTS_CNT_W(8),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o0_wo_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g0_p0_w2n_wo_icb_cmd_valid            ),
  .i0_icb_cmd_ready               (mst_g0_p0_w2n_wo_icb_cmd_ready            ),
  .i0_icb_cmd_sel                 (mst_g0_p0_w2n_wo_icb_cmd_sel             ),
  .i0_icb_cmd_read                (mst_g0_p0_w2n_wo_icb_cmd_read            ),
  .i0_icb_cmd_addr                (mst_g0_p0_w2n_wo_icb_cmd_addr [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g0_p0_w2n_wo_icb_cmd_wdata [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g0_p0_w2n_wo_icb_cmd_wmask [   7:   0]),
  .i0_icb_cmd_size                (mst_g0_p0_w2n_wo_icb_cmd_size [   2:   0]),
  .i0_icb_cmd_lock                (mst_g0_p0_w2n_wo_icb_cmd_lock            ),
  .i0_icb_cmd_excl                (mst_g0_p0_w2n_wo_icb_cmd_excl            ),
  .i0_icb_cmd_xlen                (mst_g0_p0_w2n_wo_icb_cmd_xlen [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g0_p0_w2n_wo_icb_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (mst_g0_p0_w2n_wo_icb_cmd_modes [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g0_p0_w2n_wo_icb_cmd_dmode            ),
  .i0_icb_cmd_attri               (mst_g0_p0_w2n_wo_icb_cmd_attri [   2:   0]),
  .i0_icb_cmd_beat                (mst_g0_p0_w2n_wo_icb_cmd_beat [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g0_p0_w2n_wo_icb_cmd_usr  [   2:   0]),
  .i0_icb_rsp_ready               (mst_g0_p0_w2n_wo_icb_rsp_ready            ),
  .i0_icb_rsp_valid               (mst_g0_p0_w2n_wo_icb_rsp_valid            ),
  .i0_icb_rsp_err                 (mst_g0_p0_w2n_wo_icb_rsp_err             ),
  .i0_icb_rsp_excl_ok             (mst_g0_p0_w2n_wo_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g0_p0_w2n_wo_icb_rsp_rdata [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g0_p0_w2n_wo_icb_rsp_usr  [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_0_wo_icb_cmd_valid               ),
  .o_icb_cmd_ready                (mst_grp_0_wo_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (mst_grp_0_wo_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (mst_grp_0_wo_icb_cmd_read                ),
  .o_icb_cmd_addr                 (mst_grp_0_wo_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_0_wo_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_0_wo_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_0_wo_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_0_wo_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (mst_grp_0_wo_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (mst_grp_0_wo_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_0_wo_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_0_wo_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_0_wo_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (mst_grp_0_wo_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_0_wo_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_0_wo_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_0_wo_icb_rsp_ready               ),
  .o_icb_rsp_valid                (mst_grp_0_wo_icb_rsp_valid               ),
  .o_icb_rsp_err                  (mst_grp_0_wo_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (mst_grp_0_wo_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (mst_grp_0_wo_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_0_wo_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                mst_grp_1_icb_cmd_valid       ;
  wire                mst_grp_1_icb_cmd_ready       ;
  wire                mst_grp_1_icb_cmd_sel         ;
  wire                mst_grp_1_icb_cmd_read        ;
  wire    [  31:   0] mst_grp_1_icb_cmd_addr        ;
  wire    [  63:   0] mst_grp_1_icb_cmd_wdata       ;
  wire    [   7:   0] mst_grp_1_icb_cmd_wmask       ;
  wire    [   2:   0] mst_grp_1_icb_cmd_size        ;
  wire                mst_grp_1_icb_cmd_lock        ;
  wire                mst_grp_1_icb_cmd_excl        ;
  wire    [   7:   0] mst_grp_1_icb_cmd_xlen        ;
  wire    [   1:   0] mst_grp_1_icb_cmd_xburst      ;
  wire    [   1:   0] mst_grp_1_icb_cmd_modes       ;
  wire                mst_grp_1_icb_cmd_dmode       ;
  wire    [   2:   0] mst_grp_1_icb_cmd_attri       ;
  wire    [   1:   0] mst_grp_1_icb_cmd_beat        ;
  wire    [   2:   0] mst_grp_1_icb_cmd_usr         ;
  wire                mst_grp_1_icb_rsp_ready       ;
  wire                mst_grp_1_icb_rsp_valid       ;
  wire                mst_grp_1_icb_rsp_err         ;
  wire                mst_grp_1_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_grp_1_icb_rsp_rdata       ;
  wire    [   2:   0] mst_grp_1_icb_rsp_usr         ;
                 wire                mst_g1_p0_icb_cmd_valid       ;
  wire                mst_g1_p0_icb_cmd_ready       ;
  wire                mst_g1_p0_icb_cmd_sel         ;
  wire                mst_g1_p0_icb_cmd_read        ;
  wire    [  31:   0] mst_g1_p0_icb_cmd_addr        ;
  wire    [  63:   0] mst_g1_p0_icb_cmd_wdata       ;
  wire    [   7:   0] mst_g1_p0_icb_cmd_wmask       ;
  wire    [   2:   0] mst_g1_p0_icb_cmd_size        ;
  wire                mst_g1_p0_icb_cmd_lock        ;
  wire                mst_g1_p0_icb_cmd_excl        ;
  wire    [   7:   0] mst_g1_p0_icb_cmd_xlen        ;
  wire    [   1:   0] mst_g1_p0_icb_cmd_xburst      ;
  wire    [   1:   0] mst_g1_p0_icb_cmd_modes       ;
  wire                mst_g1_p0_icb_cmd_dmode       ;
  wire    [   2:   0] mst_g1_p0_icb_cmd_attri       ;
  wire    [   1:   0] mst_g1_p0_icb_cmd_beat        ;
  wire    [   2:   0] mst_g1_p0_icb_cmd_usr         ;
  wire                mst_g1_p0_icb_rsp_ready       ;
  wire                mst_g1_p0_icb_rsp_valid       ;
  wire                mst_g1_p0_icb_rsp_err         ;
  wire                mst_g1_p0_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_g1_p0_icb_rsp_rdata       ;
  wire    [   2:   0] mst_g1_p0_icb_rsp_usr         ;
                 wire                mst_g1_p0_w2n_icb_cmd_valid   ;
  wire                mst_g1_p0_w2n_icb_cmd_ready   ;
  wire                mst_g1_p0_w2n_icb_cmd_sel     ;
  wire                mst_g1_p0_w2n_icb_cmd_read    ;
  wire    [  31:   0] mst_g1_p0_w2n_icb_cmd_addr    ;
  wire    [  63:   0] mst_g1_p0_w2n_icb_cmd_wdata   ;
  wire    [   7:   0] mst_g1_p0_w2n_icb_cmd_wmask   ;
  wire    [   2:   0] mst_g1_p0_w2n_icb_cmd_size    ;
  wire                mst_g1_p0_w2n_icb_cmd_lock    ;
  wire                mst_g1_p0_w2n_icb_cmd_excl    ;
  wire    [   7:   0] mst_g1_p0_w2n_icb_cmd_xlen    ;
  wire    [   1:   0] mst_g1_p0_w2n_icb_cmd_xburst  ;
  wire    [   1:   0] mst_g1_p0_w2n_icb_cmd_modes   ;
  wire                mst_g1_p0_w2n_icb_cmd_dmode   ;
  wire    [   2:   0] mst_g1_p0_w2n_icb_cmd_attri   ;
  wire    [   1:   0] mst_g1_p0_w2n_icb_cmd_beat    ;
  wire    [   2:   0] mst_g1_p0_w2n_icb_cmd_usr     ;
  wire                mst_g1_p0_w2n_icb_rsp_ready   ;
  wire                mst_g1_p0_w2n_icb_rsp_valid   ;
  wire                mst_g1_p0_w2n_icb_rsp_err     ;
  wire                mst_g1_p0_w2n_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g1_p0_w2n_icb_rsp_rdata   ;
  wire    [   2:   0] mst_g1_p0_w2n_icb_rsp_usr     ;
    wire udma_r_icb_bus_active;
              wire[3-1:0] mst_g1_p0_icb_cmd_usr_pre;
               assign mst_g1_p0_icb_cmd_usr_pre = 3'b0;
               assign mst_g1_p0_icb_cmd_usr = mst_g1_p0_icb_cmd_usr_pre;
    e603_subsys_gnrl_ficb_buffer # (
           .OUTS_CNT_BLOCK_THROUGH(1),
      .I_SUPPORT_RATIO(0),
      .O_SUPPORT_RATIO(0),
      .CMD_DP(2),
      .RSP_DP(2),
      .OUTS_CNT_W     (7),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .AW    (32),
      .DW    (64), 
      .CMD_CUT_READY (1),
      .RSP_CUT_READY (1),
      .RSP_ALWAYS_READY(0),
      .ACTIVE_USE_FLOP_CLEAN (1),
      .CMD_UW (1),
      .RSP_UW (1)
    )u_mst_g1_p0_icb_icb_buffer(
      .i_clk_en   (1'b1),
      .o_clk_en   (1'b1),
      .icb_buffer_active (udma_r_icb_bus_active),
      .i_icb_cmd_read(1'b1),
      .i_icb_cmd_wdata(64'b0),
      .i_icb_cmd_wmask(8'b0),
                .i_icb_cmd_usr(1'b0),
                .i_icb_rsp_usr(),
        .i_icb_cmd_valid                (udma_r_icb_cmd_valid                     ),
  .i_icb_cmd_ready                (udma_r_icb_cmd_ready                     ),
  .i_icb_cmd_sel                  (udma_r_icb_cmd_sel                       ),
  .i_icb_cmd_size                 (udma_r_icb_cmd_size           [   2:   0]),
  .i_icb_cmd_lock                 (udma_r_icb_cmd_lock                      ),
  .i_icb_cmd_excl                 (udma_r_icb_cmd_excl                      ),
  .i_icb_cmd_xlen                 (udma_r_icb_cmd_xlen           [   7:   0]),
  .i_icb_cmd_xburst               (udma_r_icb_cmd_xburst         [   1:   0]),
  .i_icb_cmd_modes                (udma_r_icb_cmd_modes          [   1:   0]),
  .i_icb_cmd_dmode                (udma_r_icb_cmd_dmode                     ),
  .i_icb_cmd_attri                (udma_r_icb_cmd_attri          [   2:   0]),
  .i_icb_cmd_beat                 (udma_r_icb_cmd_beat           [   1:   0]),
  .i_icb_rsp_ready                (udma_r_icb_rsp_ready                     ),
  .i_icb_rsp_valid                (udma_r_icb_rsp_valid                     ),
  .i_icb_rsp_err                  (udma_r_icb_rsp_err                       ),
  .i_icb_rsp_excl_ok              (udma_r_icb_rsp_excl_ok                   ),
  .i_icb_rsp_rdata                (udma_r_icb_rsp_rdata          [  63:   0]),
      .i_icb_cmd_addr(udma_r_icb_cmd_addr[32-1:0]),
                .o_icb_cmd_usr(),
                .o_icb_rsp_usr(1'b0),
        .o_icb_cmd_valid                (mst_g1_p0_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (mst_g1_p0_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (mst_g1_p0_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (mst_g1_p0_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (mst_g1_p0_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (mst_g1_p0_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (mst_g1_p0_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (mst_g1_p0_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (mst_g1_p0_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (mst_g1_p0_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (mst_g1_p0_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (mst_g1_p0_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (mst_g1_p0_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (mst_g1_p0_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (mst_g1_p0_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (mst_g1_p0_icb_cmd_beat        [   1:   0]),
  .o_icb_rsp_ready                (mst_g1_p0_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (mst_g1_p0_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (mst_g1_p0_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (mst_g1_p0_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (mst_g1_p0_icb_rsp_rdata       [  63:   0]),
      .clk  (clk),  
      .rst_n(rst_n)
    );
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g1_p0_icb_ficb_wconv(
      .i_icb_cmd_read(1'b1),
      .i_icb_cmd_wdata(64'b0),
      .i_icb_cmd_wmask(8'b0),
        .i_icb_cmd_valid                (mst_g1_p0_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (mst_g1_p0_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (mst_g1_p0_icb_cmd_sel                    ),
  .i_icb_cmd_addr                 (mst_g1_p0_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_size                 (mst_g1_p0_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (mst_g1_p0_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (mst_g1_p0_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (mst_g1_p0_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (mst_g1_p0_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (mst_g1_p0_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (mst_g1_p0_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (mst_g1_p0_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (mst_g1_p0_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (mst_g1_p0_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (mst_g1_p0_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (mst_g1_p0_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (mst_g1_p0_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (mst_g1_p0_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (mst_g1_p0_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (mst_g1_p0_icb_rsp_usr         [   2:   0]),
        .o_icb_cmd_valid                (mst_g1_p0_w2n_icb_cmd_valid              ),
  .o_icb_cmd_ready                (mst_g1_p0_w2n_icb_cmd_ready              ),
  .o_icb_cmd_sel                  (mst_g1_p0_w2n_icb_cmd_sel                ),
  .o_icb_cmd_read                 (mst_g1_p0_w2n_icb_cmd_read               ),
  .o_icb_cmd_addr                 (mst_g1_p0_w2n_icb_cmd_addr    [  31:   0]),
  .o_icb_cmd_wdata                (mst_g1_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .o_icb_cmd_wmask                (mst_g1_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .o_icb_cmd_size                 (mst_g1_p0_w2n_icb_cmd_size    [   2:   0]),
  .o_icb_cmd_lock                 (mst_g1_p0_w2n_icb_cmd_lock               ),
  .o_icb_cmd_excl                 (mst_g1_p0_w2n_icb_cmd_excl               ),
  .o_icb_cmd_xlen                 (mst_g1_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .o_icb_cmd_xburst               (mst_g1_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .o_icb_cmd_modes                (mst_g1_p0_w2n_icb_cmd_modes   [   1:   0]),
  .o_icb_cmd_dmode                (mst_g1_p0_w2n_icb_cmd_dmode              ),
  .o_icb_cmd_attri                (mst_g1_p0_w2n_icb_cmd_attri   [   2:   0]),
  .o_icb_cmd_beat                 (mst_g1_p0_w2n_icb_cmd_beat    [   1:   0]),
  .o_icb_cmd_usr                  (mst_g1_p0_w2n_icb_cmd_usr     [   2:   0]),
  .o_icb_rsp_ready                (mst_g1_p0_w2n_icb_rsp_ready              ),
  .o_icb_rsp_valid                (mst_g1_p0_w2n_icb_rsp_valid              ),
  .o_icb_rsp_err                  (mst_g1_p0_w2n_icb_rsp_err                ),
  .o_icb_rsp_excl_ok              (mst_g1_p0_w2n_icb_rsp_excl_ok            ),
  .o_icb_rsp_rdata                (mst_g1_p0_w2n_icb_rsp_rdata   [  63:   0]),
  .o_icb_rsp_usr                  (mst_g1_p0_w2n_icb_rsp_usr     [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   e603_subsys_mgrp1_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o1_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g1_p0_w2n_icb_cmd_valid              ),
  .i0_icb_cmd_ready               (mst_g1_p0_w2n_icb_cmd_ready              ),
  .i0_icb_cmd_sel                 (mst_g1_p0_w2n_icb_cmd_sel                ),
  .i0_icb_cmd_read                (mst_g1_p0_w2n_icb_cmd_read               ),
  .i0_icb_cmd_addr                (mst_g1_p0_w2n_icb_cmd_addr    [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g1_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g1_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .i0_icb_cmd_size                (mst_g1_p0_w2n_icb_cmd_size    [   2:   0]),
  .i0_icb_cmd_lock                (mst_g1_p0_w2n_icb_cmd_lock               ),
  .i0_icb_cmd_excl                (mst_g1_p0_w2n_icb_cmd_excl               ),
  .i0_icb_cmd_xlen                (mst_g1_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g1_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .i0_icb_cmd_modes               (mst_g1_p0_w2n_icb_cmd_modes   [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g1_p0_w2n_icb_cmd_dmode              ),
  .i0_icb_cmd_attri               (mst_g1_p0_w2n_icb_cmd_attri   [   2:   0]),
  .i0_icb_cmd_beat                (mst_g1_p0_w2n_icb_cmd_beat    [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g1_p0_w2n_icb_cmd_usr     [   2:   0]),
  .i0_icb_rsp_ready               (mst_g1_p0_w2n_icb_rsp_ready              ),
  .i0_icb_rsp_valid               (mst_g1_p0_w2n_icb_rsp_valid              ),
  .i0_icb_rsp_err                 (mst_g1_p0_w2n_icb_rsp_err                ),
  .i0_icb_rsp_excl_ok             (mst_g1_p0_w2n_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g1_p0_w2n_icb_rsp_rdata   [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g1_p0_w2n_icb_rsp_usr     [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_1_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (mst_grp_1_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (mst_grp_1_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (mst_grp_1_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (mst_grp_1_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_1_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_1_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_1_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_1_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (mst_grp_1_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (mst_grp_1_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_1_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_1_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_1_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (mst_grp_1_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_1_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_1_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_1_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (mst_grp_1_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (mst_grp_1_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (mst_grp_1_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (mst_grp_1_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_1_icb_rsp_usr         [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                mst_grp_2_icb_cmd_valid       ;
  wire                mst_grp_2_icb_cmd_ready       ;
  wire                mst_grp_2_icb_cmd_sel         ;
  wire                mst_grp_2_icb_cmd_read        ;
  wire    [  31:   0] mst_grp_2_icb_cmd_addr        ;
  wire    [  63:   0] mst_grp_2_icb_cmd_wdata       ;
  wire    [   7:   0] mst_grp_2_icb_cmd_wmask       ;
  wire    [   2:   0] mst_grp_2_icb_cmd_size        ;
  wire                mst_grp_2_icb_cmd_lock        ;
  wire                mst_grp_2_icb_cmd_excl        ;
  wire    [   7:   0] mst_grp_2_icb_cmd_xlen        ;
  wire    [   1:   0] mst_grp_2_icb_cmd_xburst      ;
  wire    [   1:   0] mst_grp_2_icb_cmd_modes       ;
  wire                mst_grp_2_icb_cmd_dmode       ;
  wire    [   2:   0] mst_grp_2_icb_cmd_attri       ;
  wire    [   1:   0] mst_grp_2_icb_cmd_beat        ;
  wire    [   2:   0] mst_grp_2_icb_cmd_usr         ;
  wire                mst_grp_2_icb_rsp_ready       ;
  wire                mst_grp_2_icb_rsp_valid       ;
  wire                mst_grp_2_icb_rsp_err         ;
  wire                mst_grp_2_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_grp_2_icb_rsp_rdata       ;
  wire    [   2:   0] mst_grp_2_icb_rsp_usr         ;
                 wire                mst_g2_p0_icb_cmd_valid       ;
  wire                mst_g2_p0_icb_cmd_ready       ;
  wire                mst_g2_p0_icb_cmd_sel         ;
  wire                mst_g2_p0_icb_cmd_read        ;
  wire    [  31:   0] mst_g2_p0_icb_cmd_addr        ;
  wire    [  63:   0] mst_g2_p0_icb_cmd_wdata       ;
  wire    [   7:   0] mst_g2_p0_icb_cmd_wmask       ;
  wire    [   2:   0] mst_g2_p0_icb_cmd_size        ;
  wire                mst_g2_p0_icb_cmd_lock        ;
  wire                mst_g2_p0_icb_cmd_excl        ;
  wire    [   7:   0] mst_g2_p0_icb_cmd_xlen        ;
  wire    [   1:   0] mst_g2_p0_icb_cmd_xburst      ;
  wire    [   1:   0] mst_g2_p0_icb_cmd_modes       ;
  wire                mst_g2_p0_icb_cmd_dmode       ;
  wire    [   2:   0] mst_g2_p0_icb_cmd_attri       ;
  wire    [   1:   0] mst_g2_p0_icb_cmd_beat        ;
  wire    [   2:   0] mst_g2_p0_icb_cmd_usr         ;
  wire                mst_g2_p0_icb_rsp_ready       ;
  wire                mst_g2_p0_icb_rsp_valid       ;
  wire                mst_g2_p0_icb_rsp_err         ;
  wire                mst_g2_p0_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_g2_p0_icb_rsp_rdata       ;
  wire    [   2:   0] mst_g2_p0_icb_rsp_usr         ;
                 wire                mst_g2_p0_w2n_icb_cmd_valid   ;
  wire                mst_g2_p0_w2n_icb_cmd_ready   ;
  wire                mst_g2_p0_w2n_icb_cmd_sel     ;
  wire                mst_g2_p0_w2n_icb_cmd_read    ;
  wire    [  31:   0] mst_g2_p0_w2n_icb_cmd_addr    ;
  wire    [  63:   0] mst_g2_p0_w2n_icb_cmd_wdata   ;
  wire    [   7:   0] mst_g2_p0_w2n_icb_cmd_wmask   ;
  wire    [   2:   0] mst_g2_p0_w2n_icb_cmd_size    ;
  wire                mst_g2_p0_w2n_icb_cmd_lock    ;
  wire                mst_g2_p0_w2n_icb_cmd_excl    ;
  wire    [   7:   0] mst_g2_p0_w2n_icb_cmd_xlen    ;
  wire    [   1:   0] mst_g2_p0_w2n_icb_cmd_xburst  ;
  wire    [   1:   0] mst_g2_p0_w2n_icb_cmd_modes   ;
  wire                mst_g2_p0_w2n_icb_cmd_dmode   ;
  wire    [   2:   0] mst_g2_p0_w2n_icb_cmd_attri   ;
  wire    [   1:   0] mst_g2_p0_w2n_icb_cmd_beat    ;
  wire    [   2:   0] mst_g2_p0_w2n_icb_cmd_usr     ;
  wire                mst_g2_p0_w2n_icb_rsp_ready   ;
  wire                mst_g2_p0_w2n_icb_rsp_valid   ;
  wire                mst_g2_p0_w2n_icb_rsp_err     ;
  wire                mst_g2_p0_w2n_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g2_p0_w2n_icb_rsp_rdata   ;
  wire    [   2:   0] mst_g2_p0_w2n_icb_rsp_usr     ;
    wire udma_w_icb_bus_active;
              wire[3-1:0] mst_g2_p0_icb_cmd_usr_pre;
               assign mst_g2_p0_icb_cmd_usr_pre = 3'b0;
               assign mst_g2_p0_icb_cmd_usr = mst_g2_p0_icb_cmd_usr_pre;
    e603_subsys_gnrl_ficb_buffer # (
           .OUTS_CNT_BLOCK_THROUGH(1),
      .I_SUPPORT_RATIO(0),
      .O_SUPPORT_RATIO(0),
      .CMD_DP(2),
      .RSP_DP(2),
      .OUTS_CNT_W     (7),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .AW    (32),
      .DW    (64), 
      .CMD_CUT_READY (1),
      .RSP_CUT_READY (1),
      .RSP_ALWAYS_READY(0),
      .ACTIVE_USE_FLOP_CLEAN (1),
      .CMD_UW (1),
      .RSP_UW (1)
    )u_mst_g2_p0_icb_icb_buffer(
      .i_clk_en   (1'b1),
      .o_clk_en   (1'b1),
      .icb_buffer_active (udma_w_icb_bus_active),
                .i_icb_cmd_usr(1'b0),
                .i_icb_rsp_usr(),
        .i_icb_cmd_valid                (udma_w_icb_cmd_valid                     ),
  .i_icb_cmd_ready                (udma_w_icb_cmd_ready                     ),
  .i_icb_cmd_sel                  (udma_w_icb_cmd_sel                       ),
  .i_icb_cmd_read                 (udma_w_icb_cmd_read                      ),
  .i_icb_cmd_wdata                (udma_w_icb_cmd_wdata          [  63:   0]),
  .i_icb_cmd_wmask                (udma_w_icb_cmd_wmask          [   7:   0]),
  .i_icb_cmd_size                 (udma_w_icb_cmd_size           [   2:   0]),
  .i_icb_cmd_lock                 (udma_w_icb_cmd_lock                      ),
  .i_icb_cmd_excl                 (udma_w_icb_cmd_excl                      ),
  .i_icb_cmd_xlen                 (udma_w_icb_cmd_xlen           [   7:   0]),
  .i_icb_cmd_xburst               (udma_w_icb_cmd_xburst         [   1:   0]),
  .i_icb_cmd_modes                (udma_w_icb_cmd_modes          [   1:   0]),
  .i_icb_cmd_dmode                (udma_w_icb_cmd_dmode                     ),
  .i_icb_cmd_attri                (udma_w_icb_cmd_attri          [   2:   0]),
  .i_icb_cmd_beat                 (udma_w_icb_cmd_beat           [   1:   0]),
  .i_icb_rsp_ready                (udma_w_icb_rsp_ready                     ),
  .i_icb_rsp_valid                (udma_w_icb_rsp_valid                     ),
  .i_icb_rsp_err                  (udma_w_icb_rsp_err                       ),
  .i_icb_rsp_excl_ok              (udma_w_icb_rsp_excl_ok                   ),
  .i_icb_rsp_rdata                (udma_w_icb_rsp_rdata          [  63:   0]),
      .i_icb_cmd_addr(udma_w_icb_cmd_addr[32-1:0]),
      .o_icb_rsp_rdata(64'b0),
                .o_icb_cmd_usr(),
                .o_icb_rsp_usr(1'b0),
        .o_icb_cmd_valid                (mst_g2_p0_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (mst_g2_p0_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (mst_g2_p0_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (mst_g2_p0_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (mst_g2_p0_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (mst_g2_p0_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (mst_g2_p0_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (mst_g2_p0_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (mst_g2_p0_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (mst_g2_p0_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (mst_g2_p0_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (mst_g2_p0_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (mst_g2_p0_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (mst_g2_p0_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (mst_g2_p0_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (mst_g2_p0_icb_cmd_beat        [   1:   0]),
  .o_icb_rsp_ready                (mst_g2_p0_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (mst_g2_p0_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (mst_g2_p0_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (mst_g2_p0_icb_rsp_excl_ok                ),
      .clk  (clk),  
      .rst_n(rst_n)
    );
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g2_p0_icb_ficb_wconv(
        .i_icb_cmd_valid                (mst_g2_p0_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (mst_g2_p0_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (mst_g2_p0_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (mst_g2_p0_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (mst_g2_p0_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (mst_g2_p0_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (mst_g2_p0_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (mst_g2_p0_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (mst_g2_p0_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (mst_g2_p0_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (mst_g2_p0_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (mst_g2_p0_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (mst_g2_p0_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (mst_g2_p0_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (mst_g2_p0_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (mst_g2_p0_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (mst_g2_p0_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (mst_g2_p0_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (mst_g2_p0_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (mst_g2_p0_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (mst_g2_p0_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (mst_g2_p0_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (mst_g2_p0_icb_rsp_usr         [   2:   0]),
      .o_icb_rsp_rdata(64'b0),
        .o_icb_cmd_valid                (mst_g2_p0_w2n_icb_cmd_valid              ),
  .o_icb_cmd_ready                (mst_g2_p0_w2n_icb_cmd_ready              ),
  .o_icb_cmd_sel                  (mst_g2_p0_w2n_icb_cmd_sel                ),
  .o_icb_cmd_read                 (mst_g2_p0_w2n_icb_cmd_read               ),
  .o_icb_cmd_addr                 (mst_g2_p0_w2n_icb_cmd_addr    [  31:   0]),
  .o_icb_cmd_wdata                (mst_g2_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .o_icb_cmd_wmask                (mst_g2_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .o_icb_cmd_size                 (mst_g2_p0_w2n_icb_cmd_size    [   2:   0]),
  .o_icb_cmd_lock                 (mst_g2_p0_w2n_icb_cmd_lock               ),
  .o_icb_cmd_excl                 (mst_g2_p0_w2n_icb_cmd_excl               ),
  .o_icb_cmd_xlen                 (mst_g2_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .o_icb_cmd_xburst               (mst_g2_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .o_icb_cmd_modes                (mst_g2_p0_w2n_icb_cmd_modes   [   1:   0]),
  .o_icb_cmd_dmode                (mst_g2_p0_w2n_icb_cmd_dmode              ),
  .o_icb_cmd_attri                (mst_g2_p0_w2n_icb_cmd_attri   [   2:   0]),
  .o_icb_cmd_beat                 (mst_g2_p0_w2n_icb_cmd_beat    [   1:   0]),
  .o_icb_cmd_usr                  (mst_g2_p0_w2n_icb_cmd_usr     [   2:   0]),
  .o_icb_rsp_ready                (mst_g2_p0_w2n_icb_rsp_ready              ),
  .o_icb_rsp_valid                (mst_g2_p0_w2n_icb_rsp_valid              ),
  .o_icb_rsp_err                  (mst_g2_p0_w2n_icb_rsp_err                ),
  .o_icb_rsp_excl_ok              (mst_g2_p0_w2n_icb_rsp_excl_ok            ),
  .o_icb_rsp_usr                  (mst_g2_p0_w2n_icb_rsp_usr     [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   e603_subsys_mgrp2_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o2_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g2_p0_w2n_icb_cmd_valid              ),
  .i0_icb_cmd_ready               (mst_g2_p0_w2n_icb_cmd_ready              ),
  .i0_icb_cmd_sel                 (mst_g2_p0_w2n_icb_cmd_sel                ),
  .i0_icb_cmd_read                (mst_g2_p0_w2n_icb_cmd_read               ),
  .i0_icb_cmd_addr                (mst_g2_p0_w2n_icb_cmd_addr    [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g2_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g2_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .i0_icb_cmd_size                (mst_g2_p0_w2n_icb_cmd_size    [   2:   0]),
  .i0_icb_cmd_lock                (mst_g2_p0_w2n_icb_cmd_lock               ),
  .i0_icb_cmd_excl                (mst_g2_p0_w2n_icb_cmd_excl               ),
  .i0_icb_cmd_xlen                (mst_g2_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g2_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .i0_icb_cmd_modes               (mst_g2_p0_w2n_icb_cmd_modes   [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g2_p0_w2n_icb_cmd_dmode              ),
  .i0_icb_cmd_attri               (mst_g2_p0_w2n_icb_cmd_attri   [   2:   0]),
  .i0_icb_cmd_beat                (mst_g2_p0_w2n_icb_cmd_beat    [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g2_p0_w2n_icb_cmd_usr     [   2:   0]),
  .i0_icb_rsp_ready               (mst_g2_p0_w2n_icb_rsp_ready              ),
  .i0_icb_rsp_valid               (mst_g2_p0_w2n_icb_rsp_valid              ),
  .i0_icb_rsp_err                 (mst_g2_p0_w2n_icb_rsp_err                ),
  .i0_icb_rsp_excl_ok             (mst_g2_p0_w2n_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g2_p0_w2n_icb_rsp_rdata   [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g2_p0_w2n_icb_rsp_usr     [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_2_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (mst_grp_2_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (mst_grp_2_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (mst_grp_2_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (mst_grp_2_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_2_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_2_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_2_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_2_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (mst_grp_2_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (mst_grp_2_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_2_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_2_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_2_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (mst_grp_2_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_2_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_2_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_2_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (mst_grp_2_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (mst_grp_2_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (mst_grp_2_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (mst_grp_2_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_2_icb_rsp_usr         [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                mst_grp_3_icb_cmd_valid       ;
  wire                mst_grp_3_icb_cmd_ready       ;
  wire                mst_grp_3_icb_cmd_sel         ;
  wire                mst_grp_3_icb_cmd_read        ;
  wire    [  31:   0] mst_grp_3_icb_cmd_addr        ;
  wire    [  63:   0] mst_grp_3_icb_cmd_wdata       ;
  wire    [   7:   0] mst_grp_3_icb_cmd_wmask       ;
  wire    [   2:   0] mst_grp_3_icb_cmd_size        ;
  wire                mst_grp_3_icb_cmd_lock        ;
  wire                mst_grp_3_icb_cmd_excl        ;
  wire    [   7:   0] mst_grp_3_icb_cmd_xlen        ;
  wire    [   1:   0] mst_grp_3_icb_cmd_xburst      ;
  wire    [   1:   0] mst_grp_3_icb_cmd_modes       ;
  wire                mst_grp_3_icb_cmd_dmode       ;
  wire    [   2:   0] mst_grp_3_icb_cmd_attri       ;
  wire    [   1:   0] mst_grp_3_icb_cmd_beat        ;
  wire    [   2:   0] mst_grp_3_icb_cmd_usr         ;
  wire                mst_grp_3_icb_rsp_ready       ;
  wire                mst_grp_3_icb_rsp_valid       ;
  wire                mst_grp_3_icb_rsp_err         ;
  wire                mst_grp_3_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_grp_3_icb_rsp_rdata       ;
  wire    [   2:   0] mst_grp_3_icb_rsp_usr         ;
                 wire                mst_g3_p0_icb_cmd_valid       ;
  wire                mst_g3_p0_icb_cmd_ready       ;
  wire                mst_g3_p0_icb_cmd_sel         ;
  wire                mst_g3_p0_icb_cmd_read        ;
  wire    [  31:   0] mst_g3_p0_icb_cmd_addr        ;
  wire    [  63:   0] mst_g3_p0_icb_cmd_wdata       ;
  wire    [   7:   0] mst_g3_p0_icb_cmd_wmask       ;
  wire    [   2:   0] mst_g3_p0_icb_cmd_size        ;
  wire                mst_g3_p0_icb_cmd_lock        ;
  wire                mst_g3_p0_icb_cmd_excl        ;
  wire    [   7:   0] mst_g3_p0_icb_cmd_xlen        ;
  wire    [   1:   0] mst_g3_p0_icb_cmd_xburst      ;
  wire    [   1:   0] mst_g3_p0_icb_cmd_modes       ;
  wire                mst_g3_p0_icb_cmd_dmode       ;
  wire    [   2:   0] mst_g3_p0_icb_cmd_attri       ;
  wire    [   1:   0] mst_g3_p0_icb_cmd_beat        ;
  wire    [   2:   0] mst_g3_p0_icb_cmd_usr         ;
  wire                mst_g3_p0_icb_rsp_ready       ;
  wire                mst_g3_p0_icb_rsp_valid       ;
  wire                mst_g3_p0_icb_rsp_err         ;
  wire                mst_g3_p0_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_g3_p0_icb_rsp_rdata       ;
  wire    [   2:   0] mst_g3_p0_icb_rsp_usr         ;
                 wire                mst_g3_p0_w2n_icb_cmd_valid   ;
  wire                mst_g3_p0_w2n_icb_cmd_ready   ;
  wire                mst_g3_p0_w2n_icb_cmd_sel     ;
  wire                mst_g3_p0_w2n_icb_cmd_read    ;
  wire    [  31:   0] mst_g3_p0_w2n_icb_cmd_addr    ;
  wire    [  63:   0] mst_g3_p0_w2n_icb_cmd_wdata   ;
  wire    [   7:   0] mst_g3_p0_w2n_icb_cmd_wmask   ;
  wire    [   2:   0] mst_g3_p0_w2n_icb_cmd_size    ;
  wire                mst_g3_p0_w2n_icb_cmd_lock    ;
  wire                mst_g3_p0_w2n_icb_cmd_excl    ;
  wire    [   7:   0] mst_g3_p0_w2n_icb_cmd_xlen    ;
  wire    [   1:   0] mst_g3_p0_w2n_icb_cmd_xburst  ;
  wire    [   1:   0] mst_g3_p0_w2n_icb_cmd_modes   ;
  wire                mst_g3_p0_w2n_icb_cmd_dmode   ;
  wire    [   2:   0] mst_g3_p0_w2n_icb_cmd_attri   ;
  wire    [   1:   0] mst_g3_p0_w2n_icb_cmd_beat    ;
  wire    [   2:   0] mst_g3_p0_w2n_icb_cmd_usr     ;
  wire                mst_g3_p0_w2n_icb_rsp_ready   ;
  wire                mst_g3_p0_w2n_icb_rsp_valid   ;
  wire                mst_g3_p0_w2n_icb_rsp_err     ;
  wire                mst_g3_p0_w2n_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g3_p0_w2n_icb_rsp_rdata   ;
  wire    [   2:   0] mst_g3_p0_w2n_icb_rsp_usr     ;
    wire dummy_icb_bus_active;
              wire[3-1:0] mst_g3_p0_icb_cmd_usr_pre;
               assign mst_g3_p0_icb_cmd_usr_pre = 3'b0;
               assign mst_g3_p0_icb_cmd_usr = mst_g3_p0_icb_cmd_usr_pre;
    e603_subsys_gnrl_ficb_buffer # (
           .OUTS_CNT_BLOCK_THROUGH(1),
      .I_SUPPORT_RATIO(0),
      .O_SUPPORT_RATIO(0),
      .CMD_DP(2),
      .RSP_DP(2),
      .OUTS_CNT_W     (7),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .AW    (32),
      .DW    (64), 
      .CMD_CUT_READY (1),
      .RSP_CUT_READY (1),
      .RSP_ALWAYS_READY(0),
      .ACTIVE_USE_FLOP_CLEAN (1),
      .CMD_UW (1),
      .RSP_UW (1)
    )u_mst_g3_p0_icb_icb_buffer(
      .i_clk_en   (1'b1),
      .o_clk_en   (1'b1),
      .icb_buffer_active (dummy_icb_bus_active),
                .i_icb_cmd_usr(1'b0),
                .i_icb_rsp_usr(),
        .i_icb_cmd_valid                (dummy_icb_cmd_valid                      ),
  .i_icb_cmd_ready                (dummy_icb_cmd_ready                      ),
  .i_icb_cmd_sel                  (dummy_icb_cmd_sel                        ),
  .i_icb_cmd_read                 (dummy_icb_cmd_read                       ),
  .i_icb_cmd_wdata                (dummy_icb_cmd_wdata           [  63:   0]),
  .i_icb_cmd_wmask                (dummy_icb_cmd_wmask           [   7:   0]),
  .i_icb_cmd_size                 (dummy_icb_cmd_size            [   2:   0]),
  .i_icb_cmd_lock                 (dummy_icb_cmd_lock                       ),
  .i_icb_cmd_excl                 (dummy_icb_cmd_excl                       ),
  .i_icb_cmd_xlen                 (dummy_icb_cmd_xlen            [   7:   0]),
  .i_icb_cmd_xburst               (dummy_icb_cmd_xburst          [   1:   0]),
  .i_icb_cmd_modes                (dummy_icb_cmd_modes           [   1:   0]),
  .i_icb_cmd_dmode                (dummy_icb_cmd_dmode                      ),
  .i_icb_cmd_attri                (dummy_icb_cmd_attri           [   2:   0]),
  .i_icb_cmd_beat                 (dummy_icb_cmd_beat            [   1:   0]),
  .i_icb_rsp_ready                (dummy_icb_rsp_ready                      ),
  .i_icb_rsp_valid                (dummy_icb_rsp_valid                      ),
  .i_icb_rsp_err                  (dummy_icb_rsp_err                        ),
  .i_icb_rsp_excl_ok              (dummy_icb_rsp_excl_ok                    ),
  .i_icb_rsp_rdata                (dummy_icb_rsp_rdata           [  63:   0]),
      .i_icb_cmd_addr(dummy_icb_cmd_addr[32-1:0]),
                .o_icb_cmd_usr(),
                .o_icb_rsp_usr(1'b0),
        .o_icb_cmd_valid                (mst_g3_p0_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (mst_g3_p0_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (mst_g3_p0_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (mst_g3_p0_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (mst_g3_p0_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (mst_g3_p0_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (mst_g3_p0_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (mst_g3_p0_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (mst_g3_p0_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (mst_g3_p0_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (mst_g3_p0_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (mst_g3_p0_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (mst_g3_p0_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (mst_g3_p0_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (mst_g3_p0_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (mst_g3_p0_icb_cmd_beat        [   1:   0]),
  .o_icb_rsp_ready                (mst_g3_p0_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (mst_g3_p0_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (mst_g3_p0_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (mst_g3_p0_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (mst_g3_p0_icb_rsp_rdata       [  63:   0]),
      .clk  (clk),  
      .rst_n(rst_n)
    );
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g3_p0_icb_ficb_wconv(
        .i_icb_cmd_valid                (mst_g3_p0_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (mst_g3_p0_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (mst_g3_p0_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (mst_g3_p0_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (mst_g3_p0_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (mst_g3_p0_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (mst_g3_p0_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (mst_g3_p0_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (mst_g3_p0_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (mst_g3_p0_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (mst_g3_p0_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (mst_g3_p0_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (mst_g3_p0_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (mst_g3_p0_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (mst_g3_p0_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (mst_g3_p0_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (mst_g3_p0_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (mst_g3_p0_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (mst_g3_p0_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (mst_g3_p0_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (mst_g3_p0_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (mst_g3_p0_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (mst_g3_p0_icb_rsp_usr         [   2:   0]),
        .o_icb_cmd_valid                (mst_g3_p0_w2n_icb_cmd_valid              ),
  .o_icb_cmd_ready                (mst_g3_p0_w2n_icb_cmd_ready              ),
  .o_icb_cmd_sel                  (mst_g3_p0_w2n_icb_cmd_sel                ),
  .o_icb_cmd_read                 (mst_g3_p0_w2n_icb_cmd_read               ),
  .o_icb_cmd_addr                 (mst_g3_p0_w2n_icb_cmd_addr    [  31:   0]),
  .o_icb_cmd_wdata                (mst_g3_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .o_icb_cmd_wmask                (mst_g3_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .o_icb_cmd_size                 (mst_g3_p0_w2n_icb_cmd_size    [   2:   0]),
  .o_icb_cmd_lock                 (mst_g3_p0_w2n_icb_cmd_lock               ),
  .o_icb_cmd_excl                 (mst_g3_p0_w2n_icb_cmd_excl               ),
  .o_icb_cmd_xlen                 (mst_g3_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .o_icb_cmd_xburst               (mst_g3_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .o_icb_cmd_modes                (mst_g3_p0_w2n_icb_cmd_modes   [   1:   0]),
  .o_icb_cmd_dmode                (mst_g3_p0_w2n_icb_cmd_dmode              ),
  .o_icb_cmd_attri                (mst_g3_p0_w2n_icb_cmd_attri   [   2:   0]),
  .o_icb_cmd_beat                 (mst_g3_p0_w2n_icb_cmd_beat    [   1:   0]),
  .o_icb_cmd_usr                  (mst_g3_p0_w2n_icb_cmd_usr     [   2:   0]),
  .o_icb_rsp_ready                (mst_g3_p0_w2n_icb_rsp_ready              ),
  .o_icb_rsp_valid                (mst_g3_p0_w2n_icb_rsp_valid              ),
  .o_icb_rsp_err                  (mst_g3_p0_w2n_icb_rsp_err                ),
  .o_icb_rsp_excl_ok              (mst_g3_p0_w2n_icb_rsp_excl_ok            ),
  .o_icb_rsp_rdata                (mst_g3_p0_w2n_icb_rsp_rdata   [  63:   0]),
  .o_icb_rsp_usr                  (mst_g3_p0_w2n_icb_rsp_usr     [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   e603_subsys_mgrp3_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o3_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g3_p0_w2n_icb_cmd_valid              ),
  .i0_icb_cmd_ready               (mst_g3_p0_w2n_icb_cmd_ready              ),
  .i0_icb_cmd_sel                 (mst_g3_p0_w2n_icb_cmd_sel                ),
  .i0_icb_cmd_read                (mst_g3_p0_w2n_icb_cmd_read               ),
  .i0_icb_cmd_addr                (mst_g3_p0_w2n_icb_cmd_addr    [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g3_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g3_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .i0_icb_cmd_size                (mst_g3_p0_w2n_icb_cmd_size    [   2:   0]),
  .i0_icb_cmd_lock                (mst_g3_p0_w2n_icb_cmd_lock               ),
  .i0_icb_cmd_excl                (mst_g3_p0_w2n_icb_cmd_excl               ),
  .i0_icb_cmd_xlen                (mst_g3_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g3_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .i0_icb_cmd_modes               (mst_g3_p0_w2n_icb_cmd_modes   [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g3_p0_w2n_icb_cmd_dmode              ),
  .i0_icb_cmd_attri               (mst_g3_p0_w2n_icb_cmd_attri   [   2:   0]),
  .i0_icb_cmd_beat                (mst_g3_p0_w2n_icb_cmd_beat    [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g3_p0_w2n_icb_cmd_usr     [   2:   0]),
  .i0_icb_rsp_ready               (mst_g3_p0_w2n_icb_rsp_ready              ),
  .i0_icb_rsp_valid               (mst_g3_p0_w2n_icb_rsp_valid              ),
  .i0_icb_rsp_err                 (mst_g3_p0_w2n_icb_rsp_err                ),
  .i0_icb_rsp_excl_ok             (mst_g3_p0_w2n_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g3_p0_w2n_icb_rsp_rdata   [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g3_p0_w2n_icb_rsp_usr     [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_3_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (mst_grp_3_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (mst_grp_3_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (mst_grp_3_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (mst_grp_3_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_3_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_3_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_3_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_3_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (mst_grp_3_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (mst_grp_3_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_3_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_3_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_3_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (mst_grp_3_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_3_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_3_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_3_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (mst_grp_3_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (mst_grp_3_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (mst_grp_3_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (mst_grp_3_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_3_icb_rsp_usr         [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                mst_grp_4_ro_icb_cmd_valid    ;
  wire                mst_grp_4_ro_icb_cmd_ready    ;
  wire                mst_grp_4_ro_icb_cmd_sel      ;
  wire                mst_grp_4_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_4_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_4_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_4_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_4_ro_icb_cmd_size     ;
  wire                mst_grp_4_ro_icb_cmd_lock     ;
  wire                mst_grp_4_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_4_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_4_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_4_ro_icb_cmd_modes    ;
  wire                mst_grp_4_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_4_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_4_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_4_ro_icb_cmd_usr      ;
  wire                mst_grp_4_ro_icb_rsp_ready    ;
  wire                mst_grp_4_ro_icb_rsp_valid    ;
  wire                mst_grp_4_ro_icb_rsp_err      ;
  wire                mst_grp_4_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_4_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_4_ro_icb_rsp_usr      ;
      wire                mst_grp_4_wo_icb_cmd_valid    ;
  wire                mst_grp_4_wo_icb_cmd_ready    ;
  wire                mst_grp_4_wo_icb_cmd_sel      ;
  wire                mst_grp_4_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_4_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_4_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_4_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_4_wo_icb_cmd_size     ;
  wire                mst_grp_4_wo_icb_cmd_lock     ;
  wire                mst_grp_4_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_4_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_4_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_4_wo_icb_cmd_modes    ;
  wire                mst_grp_4_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_4_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_4_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_4_wo_icb_cmd_usr      ;
  wire                mst_grp_4_wo_icb_rsp_ready    ;
  wire                mst_grp_4_wo_icb_rsp_valid    ;
  wire                mst_grp_4_wo_icb_rsp_err      ;
  wire                mst_grp_4_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_4_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_4_wo_icb_rsp_usr      ;
                 wire                mst_g4_p0_icb_cmd_valid       ;
  wire                mst_g4_p0_icb_cmd_ready       ;
  wire                mst_g4_p0_icb_cmd_sel         ;
  wire                mst_g4_p0_icb_cmd_read        ;
  wire    [  31:   0] mst_g4_p0_icb_cmd_addr        ;
  wire    [  63:   0] mst_g4_p0_icb_cmd_wdata       ;
  wire    [   7:   0] mst_g4_p0_icb_cmd_wmask       ;
  wire    [   2:   0] mst_g4_p0_icb_cmd_size        ;
  wire                mst_g4_p0_icb_cmd_lock        ;
  wire                mst_g4_p0_icb_cmd_excl        ;
  wire    [   7:   0] mst_g4_p0_icb_cmd_xlen        ;
  wire    [   1:   0] mst_g4_p0_icb_cmd_xburst      ;
  wire    [   1:   0] mst_g4_p0_icb_cmd_modes       ;
  wire                mst_g4_p0_icb_cmd_dmode       ;
  wire    [   2:   0] mst_g4_p0_icb_cmd_attri       ;
  wire    [   1:   0] mst_g4_p0_icb_cmd_beat        ;
  wire    [   2:   0] mst_g4_p0_icb_cmd_usr         ;
  wire                mst_g4_p0_icb_rsp_ready       ;
  wire                mst_g4_p0_icb_rsp_valid       ;
  wire                mst_g4_p0_icb_rsp_err         ;
  wire                mst_g4_p0_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_g4_p0_icb_rsp_rdata       ;
  wire    [   2:   0] mst_g4_p0_icb_rsp_usr         ;
                wire [3-1:0] mst_g4_p0_icb_cmd_id;
                wire [3-1:0] mst_g4_p0_icb_rsp_id;
                wire                  mst_g4_p0_icb_rsp_last;
                 wire                mst_g4_p0_w2n_ro_icb_cmd_valid ;
  wire                mst_g4_p0_w2n_ro_icb_cmd_ready ;
  wire                mst_g4_p0_w2n_ro_icb_cmd_sel  ;
  wire                mst_g4_p0_w2n_ro_icb_cmd_read ;
  wire    [  31:   0] mst_g4_p0_w2n_ro_icb_cmd_addr ;
  wire    [  63:   0] mst_g4_p0_w2n_ro_icb_cmd_wdata ;
  wire    [   7:   0] mst_g4_p0_w2n_ro_icb_cmd_wmask ;
  wire    [   2:   0] mst_g4_p0_w2n_ro_icb_cmd_size ;
  wire                mst_g4_p0_w2n_ro_icb_cmd_lock ;
  wire                mst_g4_p0_w2n_ro_icb_cmd_excl ;
  wire    [   7:   0] mst_g4_p0_w2n_ro_icb_cmd_xlen ;
  wire    [   1:   0] mst_g4_p0_w2n_ro_icb_cmd_xburst ;
  wire    [   1:   0] mst_g4_p0_w2n_ro_icb_cmd_modes ;
  wire                mst_g4_p0_w2n_ro_icb_cmd_dmode ;
  wire    [   2:   0] mst_g4_p0_w2n_ro_icb_cmd_attri ;
  wire    [   1:   0] mst_g4_p0_w2n_ro_icb_cmd_beat ;
  wire    [   2:   0] mst_g4_p0_w2n_ro_icb_cmd_usr  ;
  wire                mst_g4_p0_w2n_ro_icb_rsp_ready ;
  wire                mst_g4_p0_w2n_ro_icb_rsp_valid ;
  wire                mst_g4_p0_w2n_ro_icb_rsp_err  ;
  wire                mst_g4_p0_w2n_ro_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g4_p0_w2n_ro_icb_rsp_rdata ;
  wire    [   2:   0] mst_g4_p0_w2n_ro_icb_rsp_usr  ;
                 wire                mst_g4_p0_w2n_wo_icb_cmd_valid ;
  wire                mst_g4_p0_w2n_wo_icb_cmd_ready ;
  wire                mst_g4_p0_w2n_wo_icb_cmd_sel  ;
  wire                mst_g4_p0_w2n_wo_icb_cmd_read ;
  wire    [  31:   0] mst_g4_p0_w2n_wo_icb_cmd_addr ;
  wire    [  63:   0] mst_g4_p0_w2n_wo_icb_cmd_wdata ;
  wire    [   7:   0] mst_g4_p0_w2n_wo_icb_cmd_wmask ;
  wire    [   2:   0] mst_g4_p0_w2n_wo_icb_cmd_size ;
  wire                mst_g4_p0_w2n_wo_icb_cmd_lock ;
  wire                mst_g4_p0_w2n_wo_icb_cmd_excl ;
  wire    [   7:   0] mst_g4_p0_w2n_wo_icb_cmd_xlen ;
  wire    [   1:   0] mst_g4_p0_w2n_wo_icb_cmd_xburst ;
  wire    [   1:   0] mst_g4_p0_w2n_wo_icb_cmd_modes ;
  wire                mst_g4_p0_w2n_wo_icb_cmd_dmode ;
  wire    [   2:   0] mst_g4_p0_w2n_wo_icb_cmd_attri ;
  wire    [   1:   0] mst_g4_p0_w2n_wo_icb_cmd_beat ;
  wire    [   2:   0] mst_g4_p0_w2n_wo_icb_cmd_usr  ;
  wire                mst_g4_p0_w2n_wo_icb_rsp_ready ;
  wire                mst_g4_p0_w2n_wo_icb_rsp_valid ;
  wire                mst_g4_p0_w2n_wo_icb_rsp_err  ;
  wire                mst_g4_p0_w2n_wo_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g4_p0_w2n_wo_icb_rsp_rdata ;
  wire    [   2:   0] mst_g4_p0_w2n_wo_icb_rsp_usr  ;
    wire dummy_axi_bus_active;
                 wire                mst_g4_p0_ro_icb_cmd_valid    ;
  wire                mst_g4_p0_ro_icb_cmd_ready    ;
  wire                mst_g4_p0_ro_icb_cmd_sel      ;
  wire                mst_g4_p0_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_g4_p0_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_g4_p0_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_g4_p0_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_g4_p0_ro_icb_cmd_size     ;
  wire                mst_g4_p0_ro_icb_cmd_lock     ;
  wire                mst_g4_p0_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_g4_p0_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_g4_p0_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_g4_p0_ro_icb_cmd_modes    ;
  wire                mst_g4_p0_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_g4_p0_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_g4_p0_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_g4_p0_ro_icb_cmd_usr      ;
  wire                mst_g4_p0_ro_icb_rsp_ready    ;
  wire                mst_g4_p0_ro_icb_rsp_valid    ;
  wire                mst_g4_p0_ro_icb_rsp_err      ;
  wire                mst_g4_p0_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_g4_p0_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_g4_p0_ro_icb_rsp_usr      ;
                    wire [3-1:0] mst_g4_p0_ro_icb_cmd_id;
                    wire [3-1:0] mst_g4_p0_ro_icb_rsp_id;
                    wire                  mst_g4_p0_ro_icb_rsp_last;
    wire mst_g4_p0_ro_icb_bus_active;
                              wire[3-1:0] mst_g4_p0_ro_icb_cmd_usr_pre;
               assign mst_g4_p0_ro_icb_cmd_usr = mst_g4_p0_ro_icb_cmd_usr_pre;
  e603_subsys_gnrl_axi2ficb_read_id # (
      .ALLOW_FIX_BURST(1),
      .ID_W(3),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .RATIO_FIFO_DP(2),
      .AW(32),
      .DW(64), 
      .MW(64/8), 
      .FIFO_OUTS_NUM (64),
      .USR_W (3)
    )u_dummy_axi_axi2ficb_read(
  .reset_flag_r  (1'b0),
  .axi_bus_clk_en(1'b1),
  .icb_clk_en(1'b1),
      .axi_arvalid                    (dummy_axi_arvalid                        ),
  .axi_arready                    (dummy_axi_arready                        ),
  .axi_arlen                      (dummy_axi_arlen               [   7:   0]),
  .axi_arsize                     (dummy_axi_arsize              [   2:   0]),
  .axi_arburst                    (dummy_axi_arburst             [   1:   0]),
  .axi_arlock                     (dummy_axi_arlock                         ),
  .axi_arcache                    (dummy_axi_arcache             [   3:   0]),
  .axi_arprot                     (dummy_axi_arprot              [   2:   0]),
  .axi_rready                     (dummy_axi_rready                         ),
  .axi_rvalid                     (dummy_axi_rvalid                         ),
  .axi_rdata                      (dummy_axi_rdata               [  63:   0]),
  .axi_rresp                      (dummy_axi_rresp               [   1:   0]),
  .axi_rlast                      (dummy_axi_rlast                          ),
      .axi_araddr(dummy_axi_araddr[32-1:0]),
      .axi_aruser(3'b0),
      .axi_ruser(),
      .axi_arid(dummy_axi_arid),
      .axi_rid (dummy_axi_rid ),
        .icb_rcmd_valid                 (mst_g4_p0_ro_icb_cmd_valid               ),
  .icb_rcmd_ready                 (mst_g4_p0_ro_icb_cmd_ready               ),
  .icb_rcmd_sel                   (mst_g4_p0_ro_icb_cmd_sel                 ),
  .icb_rcmd_read                  (mst_g4_p0_ro_icb_cmd_read                ),
  .icb_rcmd_addr                  (mst_g4_p0_ro_icb_cmd_addr     [  31:   0]),
  .icb_rcmd_wdata                 (mst_g4_p0_ro_icb_cmd_wdata    [  63:   0]),
  .icb_rcmd_wmask                 (mst_g4_p0_ro_icb_cmd_wmask    [   7:   0]),
  .icb_rcmd_size                  (mst_g4_p0_ro_icb_cmd_size     [   2:   0]),
  .icb_rcmd_excl                  (mst_g4_p0_ro_icb_cmd_excl                ),
  .icb_rcmd_xlen                  (mst_g4_p0_ro_icb_cmd_xlen     [   7:   0]),
  .icb_rcmd_xburst                (mst_g4_p0_ro_icb_cmd_xburst   [   1:   0]),
  .icb_rcmd_modes                 (mst_g4_p0_ro_icb_cmd_modes    [   1:   0]),
  .icb_rcmd_dmode                 (mst_g4_p0_ro_icb_cmd_dmode               ),
  .icb_rcmd_attri                 (mst_g4_p0_ro_icb_cmd_attri    [   2:   0]),
  .icb_rcmd_beat                  (mst_g4_p0_ro_icb_cmd_beat     [   1:   0]),
  .icb_rrsp_ready                 (mst_g4_p0_ro_icb_rsp_ready               ),
  .icb_rrsp_valid                 (mst_g4_p0_ro_icb_rsp_valid               ),
  .icb_rrsp_err                   (mst_g4_p0_ro_icb_rsp_err                 ),
  .icb_rrsp_excl_ok               (mst_g4_p0_ro_icb_rsp_excl_ok             ),
  .icb_rrsp_rdata                 (mst_g4_p0_ro_icb_rsp_rdata    [  63:   0]),
      .icb_rcmd_usr(mst_g4_p0_ro_icb_cmd_usr_pre),
      .icb_rrsp_usr(mst_g4_p0_ro_icb_rsp_usr[3-1:0]),
      .icb_rcmd_id(mst_g4_p0_ro_icb_cmd_id),
      .icb_rrsp_id(mst_g4_p0_ro_icb_rsp_id),
      .icb_rrsp_last(mst_g4_p0_ro_icb_rsp_last),
      .axi2icb_read_active (mst_g4_p0_ro_icb_bus_active),
      .clk  (clk_fab),  
      .rst_n(rst_n)
    );
    assign mst_g4_p0_ro_icb_cmd_lock = 1'b0;
                 wire                mst_g4_p0_wo_icb_cmd_valid    ;
  wire                mst_g4_p0_wo_icb_cmd_ready    ;
  wire                mst_g4_p0_wo_icb_cmd_sel      ;
  wire                mst_g4_p0_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_g4_p0_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_g4_p0_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_g4_p0_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_g4_p0_wo_icb_cmd_size     ;
  wire                mst_g4_p0_wo_icb_cmd_lock     ;
  wire                mst_g4_p0_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_g4_p0_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_g4_p0_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_g4_p0_wo_icb_cmd_modes    ;
  wire                mst_g4_p0_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_g4_p0_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_g4_p0_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_g4_p0_wo_icb_cmd_usr      ;
  wire                mst_g4_p0_wo_icb_rsp_ready    ;
  wire                mst_g4_p0_wo_icb_rsp_valid    ;
  wire                mst_g4_p0_wo_icb_rsp_err      ;
  wire                mst_g4_p0_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_g4_p0_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_g4_p0_wo_icb_rsp_usr      ;
                    wire [3-1:0] mst_g4_p0_wo_icb_cmd_id;
                    wire [3-1:0] mst_g4_p0_wo_icb_rsp_id;
                    wire                  mst_g4_p0_wo_icb_rsp_last;
    wire mst_g4_p0_wo_icb_bus_active;
                              wire[3-1:0] mst_g4_p0_wo_icb_cmd_usr_pre;
               assign mst_g4_p0_wo_icb_cmd_usr = mst_g4_p0_wo_icb_cmd_usr_pre;
  e603_subsys_gnrl_axi2ficb_write_id # (
      .ALLOW_FIX_BURST(1),
      .ID_W(3),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .RATIO_FIFO_DP(2),
      .AW(32),
      .DW(64), 
      .MW(64/8), 
      .FIFO_OUTS_NUM (64),
      .USR_W (3)
    )u_mst_g4_p0_wo_icb_axi2ficb_write(
  .reset_flag_r  (1'b0),
  .axi_bus_clk_en(1'b1),
  .icb_clk_en(1'b1),
      .axi_awvalid                    (dummy_axi_awvalid                        ),
  .axi_awready                    (dummy_axi_awready                        ),
  .axi_awlen                      (dummy_axi_awlen               [   7:   0]),
  .axi_awsize                     (dummy_axi_awsize              [   2:   0]),
  .axi_awburst                    (dummy_axi_awburst             [   1:   0]),
  .axi_awlock                     (dummy_axi_awlock                         ),
  .axi_awcache                    (dummy_axi_awcache             [   3:   0]),
  .axi_awprot                     (dummy_axi_awprot              [   2:   0]),
  .axi_bready                     (dummy_axi_bready                         ),
  .axi_bvalid                     (dummy_axi_bvalid                         ),
  .axi_bresp                      (dummy_axi_bresp               [   1:   0]),
  .axi_wready                     (dummy_axi_wready                         ),
  .axi_wvalid                     (dummy_axi_wvalid                         ),
  .axi_wdata                      (dummy_axi_wdata               [  63:   0]),
  .axi_wstrb                      (dummy_axi_wstrb               [   7:   0]),
  .axi_wlast                      (dummy_axi_wlast                          ),
      .axi_awaddr(dummy_axi_awaddr[32-1:0]),
      .axi_awuser(3'b0),
      .axi_buser(),
      .axi_awid(dummy_axi_awid),
      .axi_bid (dummy_axi_bid ),
        .icb_wcmd_valid                 (mst_g4_p0_wo_icb_cmd_valid               ),
  .icb_wcmd_ready                 (mst_g4_p0_wo_icb_cmd_ready               ),
  .icb_wcmd_sel                   (mst_g4_p0_wo_icb_cmd_sel                 ),
  .icb_wcmd_read                  (mst_g4_p0_wo_icb_cmd_read                ),
  .icb_wcmd_addr                  (mst_g4_p0_wo_icb_cmd_addr     [  31:   0]),
  .icb_wcmd_wdata                 (mst_g4_p0_wo_icb_cmd_wdata    [  63:   0]),
  .icb_wcmd_wmask                 (mst_g4_p0_wo_icb_cmd_wmask    [   7:   0]),
  .icb_wcmd_size                  (mst_g4_p0_wo_icb_cmd_size     [   2:   0]),
  .icb_wcmd_lock                  (mst_g4_p0_wo_icb_cmd_lock                ),
  .icb_wcmd_excl                  (mst_g4_p0_wo_icb_cmd_excl                ),
  .icb_wcmd_xlen                  (mst_g4_p0_wo_icb_cmd_xlen     [   7:   0]),
  .icb_wcmd_xburst                (mst_g4_p0_wo_icb_cmd_xburst   [   1:   0]),
  .icb_wcmd_modes                 (mst_g4_p0_wo_icb_cmd_modes    [   1:   0]),
  .icb_wcmd_dmode                 (mst_g4_p0_wo_icb_cmd_dmode               ),
  .icb_wcmd_attri                 (mst_g4_p0_wo_icb_cmd_attri    [   2:   0]),
  .icb_wcmd_beat                  (mst_g4_p0_wo_icb_cmd_beat     [   1:   0]),
  .icb_wrsp_ready                 (mst_g4_p0_wo_icb_rsp_ready               ),
  .icb_wrsp_valid                 (mst_g4_p0_wo_icb_rsp_valid               ),
  .icb_wrsp_err                   (mst_g4_p0_wo_icb_rsp_err                 ),
  .icb_wrsp_excl_ok               (mst_g4_p0_wo_icb_rsp_excl_ok             ),
      .icb_wcmd_usr(mst_g4_p0_wo_icb_cmd_usr_pre),
      .icb_wrsp_usr(mst_g4_p0_wo_icb_rsp_usr[3-1:0]),
      .icb_wcmd_id(mst_g4_p0_wo_icb_cmd_id),
      .icb_wrsp_id(mst_g4_p0_wo_icb_rsp_id),
      .axi2icb_write_active (mst_g4_p0_wo_icb_bus_active),
      .clk  (clk_fab),  
      .rst_n(rst_n)
    );
   assign dummy_axi_bus_active = 1'b0
                     | mst_g4_p0_ro_icb_bus_active
                     | mst_g4_p0_wo_icb_bus_active
                 ;
   wire mst_g4_p0_ro_icb_id_gen_ready;
   wire [1:0] mst_g4_p0_ro_icb_cmd_beat_raw;
   wire [7:0] mst_g4_p0_ro_icb_cmd_xlen_raw;
   e603_subsys_gnrl_ficb_id_gen # (
     .OUTS_FIFO_DP (64+1),
     .ID_W         (3)
   ) u_mst_g4_p0_ro_icb_ficb_id_gen(
     .i_icb_cmd_valid(mst_g4_p0_ro_icb_cmd_valid), 
     .i_icb_cmd_ready(mst_g4_p0_ro_icb_cmd_ready), 
     .i_icb_cmd_id   (mst_g4_p0_ro_icb_cmd_id),
     .i_icb_cmd_xburst (mst_g4_p0_ro_icb_cmd_xburst),
     .i_icb_cmd_beat   (mst_g4_p0_ro_icb_cmd_beat),
     .i_icb_cmd_xlen   (mst_g4_p0_ro_icb_cmd_xlen),
     .i_icb_cmd_size   (mst_g4_p0_ro_icb_cmd_size),
     .o_icb_cmd_beat   (mst_g4_p0_ro_icb_cmd_beat_raw),
     .o_icb_cmd_xlen   (mst_g4_p0_ro_icb_cmd_xlen_raw),
     .ficb_id_gen_ready (mst_g4_p0_ro_icb_id_gen_ready),
     .i_icb_rsp_valid(mst_g4_p0_ro_icb_rsp_valid), 
     .i_icb_rsp_ready(mst_g4_p0_ro_icb_rsp_ready), 
     .i_icb_rsp_id   (mst_g4_p0_ro_icb_rsp_id),
     .i_icb_rsp_last   (mst_g4_p0_ro_icb_rsp_last),
    .clk  (clk_fab),  
    .rst_n(rst_n)
     );
    wire mst_g4_p0_ro_icb_cmd_valid_raw;
    wire mst_g4_p0_ro_icb_cmd_ready_raw;
    assign mst_g4_p0_ro_icb_cmd_valid_raw = (mst_g4_p0_ro_icb_id_gen_ready) & mst_g4_p0_ro_icb_cmd_valid;
    assign mst_g4_p0_ro_icb_cmd_ready     = (mst_g4_p0_ro_icb_id_gen_ready) & mst_g4_p0_ro_icb_cmd_ready_raw;
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g4_p0_ro_icb_ficb_wconv(
      .i_icb_cmd_read(1'b1),
                .i_icb_cmd_wdata (64'b0),
                .i_icb_cmd_wmask (8'b0),
                .i_icb_cmd_valid(mst_g4_p0_ro_icb_cmd_valid_raw),
                .i_icb_cmd_ready(mst_g4_p0_ro_icb_cmd_ready_raw),
                .i_icb_cmd_beat (mst_g4_p0_ro_icb_cmd_beat_raw),
                .i_icb_cmd_xlen (mst_g4_p0_ro_icb_cmd_xlen_raw),
        .i_icb_cmd_sel                  (mst_g4_p0_ro_icb_cmd_sel                 ),
  .i_icb_cmd_addr                 (mst_g4_p0_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_size                 (mst_g4_p0_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_g4_p0_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_g4_p0_ro_icb_cmd_excl                ),
  .i_icb_cmd_xburst               (mst_g4_p0_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_g4_p0_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_g4_p0_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_g4_p0_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_usr                  (mst_g4_p0_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_g4_p0_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_g4_p0_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_g4_p0_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_g4_p0_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_g4_p0_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_g4_p0_ro_icb_rsp_usr      [   2:   0]),
        .o_icb_cmd_valid                (mst_g4_p0_w2n_ro_icb_cmd_valid            ),
  .o_icb_cmd_ready                (mst_g4_p0_w2n_ro_icb_cmd_ready            ),
  .o_icb_cmd_sel                  (mst_g4_p0_w2n_ro_icb_cmd_sel             ),
  .o_icb_cmd_read                 (mst_g4_p0_w2n_ro_icb_cmd_read            ),
  .o_icb_cmd_addr                 (mst_g4_p0_w2n_ro_icb_cmd_addr [  31:   0]),
  .o_icb_cmd_wdata                (mst_g4_p0_w2n_ro_icb_cmd_wdata [  63:   0]),
  .o_icb_cmd_wmask                (mst_g4_p0_w2n_ro_icb_cmd_wmask [   7:   0]),
  .o_icb_cmd_size                 (mst_g4_p0_w2n_ro_icb_cmd_size [   2:   0]),
  .o_icb_cmd_lock                 (mst_g4_p0_w2n_ro_icb_cmd_lock            ),
  .o_icb_cmd_excl                 (mst_g4_p0_w2n_ro_icb_cmd_excl            ),
  .o_icb_cmd_xlen                 (mst_g4_p0_w2n_ro_icb_cmd_xlen [   7:   0]),
  .o_icb_cmd_xburst               (mst_g4_p0_w2n_ro_icb_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (mst_g4_p0_w2n_ro_icb_cmd_modes [   1:   0]),
  .o_icb_cmd_dmode                (mst_g4_p0_w2n_ro_icb_cmd_dmode            ),
  .o_icb_cmd_attri                (mst_g4_p0_w2n_ro_icb_cmd_attri [   2:   0]),
  .o_icb_cmd_beat                 (mst_g4_p0_w2n_ro_icb_cmd_beat [   1:   0]),
  .o_icb_cmd_usr                  (mst_g4_p0_w2n_ro_icb_cmd_usr  [   2:   0]),
  .o_icb_rsp_ready                (mst_g4_p0_w2n_ro_icb_rsp_ready            ),
  .o_icb_rsp_valid                (mst_g4_p0_w2n_ro_icb_rsp_valid            ),
  .o_icb_rsp_err                  (mst_g4_p0_w2n_ro_icb_rsp_err             ),
  .o_icb_rsp_excl_ok              (mst_g4_p0_w2n_ro_icb_rsp_excl_ok            ),
  .o_icb_rsp_rdata                (mst_g4_p0_w2n_ro_icb_rsp_rdata [  63:   0]),
  .o_icb_rsp_usr                  (mst_g4_p0_w2n_ro_icb_rsp_usr  [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   wire mst_g4_p0_wo_icb_id_gen_ready;
   wire [1:0] mst_g4_p0_wo_icb_cmd_beat_raw;
   wire [7:0] mst_g4_p0_wo_icb_cmd_xlen_raw;
   e603_subsys_gnrl_ficb_id_gen # (
     .OUTS_FIFO_DP (64+1),
     .ID_W         (3)
   ) u_mst_g4_p0_wo_icb_ficb_id_gen(
     .i_icb_cmd_valid(mst_g4_p0_wo_icb_cmd_valid), 
     .i_icb_cmd_ready(mst_g4_p0_wo_icb_cmd_ready), 
     .i_icb_cmd_id   (mst_g4_p0_wo_icb_cmd_id),
     .i_icb_cmd_xburst (mst_g4_p0_wo_icb_cmd_xburst),
     .i_icb_cmd_beat   (mst_g4_p0_wo_icb_cmd_beat),
     .i_icb_cmd_xlen   (mst_g4_p0_wo_icb_cmd_xlen),
     .i_icb_cmd_size   (mst_g4_p0_wo_icb_cmd_size),
     .o_icb_cmd_beat   (mst_g4_p0_wo_icb_cmd_beat_raw),
     .o_icb_cmd_xlen   (mst_g4_p0_wo_icb_cmd_xlen_raw),
     .ficb_id_gen_ready (mst_g4_p0_wo_icb_id_gen_ready),
     .i_icb_rsp_valid(mst_g4_p0_wo_icb_rsp_valid), 
     .i_icb_rsp_ready(mst_g4_p0_wo_icb_rsp_ready), 
     .i_icb_rsp_id   (mst_g4_p0_wo_icb_rsp_id),
     .i_icb_rsp_last   (mst_g4_p0_wo_icb_rsp_last),
    .clk  (clk_fab),  
    .rst_n(rst_n)
     );
    wire mst_g4_p0_wo_icb_cmd_valid_raw;
    wire mst_g4_p0_wo_icb_cmd_ready_raw;
    assign mst_g4_p0_wo_icb_cmd_valid_raw = (mst_g4_p0_wo_icb_id_gen_ready) & mst_g4_p0_wo_icb_cmd_valid;
    assign mst_g4_p0_wo_icb_cmd_ready     = (mst_g4_p0_wo_icb_id_gen_ready) & mst_g4_p0_wo_icb_cmd_ready_raw;
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g4_p0_wo_icb_ficb_wconv(
                .i_icb_cmd_valid(mst_g4_p0_wo_icb_cmd_valid_raw),
                .i_icb_cmd_ready(mst_g4_p0_wo_icb_cmd_ready_raw),
                .i_icb_cmd_xlen (mst_g4_p0_wo_icb_cmd_xlen_raw),
                .i_icb_cmd_beat (mst_g4_p0_wo_icb_cmd_beat_raw),
        .i_icb_cmd_sel                  (mst_g4_p0_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_g4_p0_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_g4_p0_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_g4_p0_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_g4_p0_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_g4_p0_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_g4_p0_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_g4_p0_wo_icb_cmd_excl                ),
  .i_icb_cmd_xburst               (mst_g4_p0_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_g4_p0_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_g4_p0_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_g4_p0_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_usr                  (mst_g4_p0_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_g4_p0_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_g4_p0_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_g4_p0_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_g4_p0_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_g4_p0_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_g4_p0_wo_icb_rsp_usr      [   2:   0]),
                .o_icb_rsp_rdata (64'b0),
        .o_icb_cmd_valid                (mst_g4_p0_w2n_wo_icb_cmd_valid            ),
  .o_icb_cmd_ready                (mst_g4_p0_w2n_wo_icb_cmd_ready            ),
  .o_icb_cmd_sel                  (mst_g4_p0_w2n_wo_icb_cmd_sel             ),
  .o_icb_cmd_read                 (mst_g4_p0_w2n_wo_icb_cmd_read            ),
  .o_icb_cmd_addr                 (mst_g4_p0_w2n_wo_icb_cmd_addr [  31:   0]),
  .o_icb_cmd_wdata                (mst_g4_p0_w2n_wo_icb_cmd_wdata [  63:   0]),
  .o_icb_cmd_wmask                (mst_g4_p0_w2n_wo_icb_cmd_wmask [   7:   0]),
  .o_icb_cmd_size                 (mst_g4_p0_w2n_wo_icb_cmd_size [   2:   0]),
  .o_icb_cmd_lock                 (mst_g4_p0_w2n_wo_icb_cmd_lock            ),
  .o_icb_cmd_excl                 (mst_g4_p0_w2n_wo_icb_cmd_excl            ),
  .o_icb_cmd_xlen                 (mst_g4_p0_w2n_wo_icb_cmd_xlen [   7:   0]),
  .o_icb_cmd_xburst               (mst_g4_p0_w2n_wo_icb_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (mst_g4_p0_w2n_wo_icb_cmd_modes [   1:   0]),
  .o_icb_cmd_dmode                (mst_g4_p0_w2n_wo_icb_cmd_dmode            ),
  .o_icb_cmd_attri                (mst_g4_p0_w2n_wo_icb_cmd_attri [   2:   0]),
  .o_icb_cmd_beat                 (mst_g4_p0_w2n_wo_icb_cmd_beat [   1:   0]),
  .o_icb_cmd_usr                  (mst_g4_p0_w2n_wo_icb_cmd_usr  [   2:   0]),
  .o_icb_rsp_ready                (mst_g4_p0_w2n_wo_icb_rsp_ready            ),
  .o_icb_rsp_valid                (mst_g4_p0_w2n_wo_icb_rsp_valid            ),
  .o_icb_rsp_err                  (mst_g4_p0_w2n_wo_icb_rsp_err             ),
  .o_icb_rsp_excl_ok              (mst_g4_p0_w2n_wo_icb_rsp_excl_ok            ),
  .o_icb_rsp_usr                  (mst_g4_p0_w2n_wo_icb_rsp_usr  [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   e603_subsys_mgrp4_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o4_ro_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g4_p0_w2n_ro_icb_cmd_valid            ),
  .i0_icb_cmd_ready               (mst_g4_p0_w2n_ro_icb_cmd_ready            ),
  .i0_icb_cmd_sel                 (mst_g4_p0_w2n_ro_icb_cmd_sel             ),
  .i0_icb_cmd_read                (mst_g4_p0_w2n_ro_icb_cmd_read            ),
  .i0_icb_cmd_addr                (mst_g4_p0_w2n_ro_icb_cmd_addr [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g4_p0_w2n_ro_icb_cmd_wdata [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g4_p0_w2n_ro_icb_cmd_wmask [   7:   0]),
  .i0_icb_cmd_size                (mst_g4_p0_w2n_ro_icb_cmd_size [   2:   0]),
  .i0_icb_cmd_lock                (mst_g4_p0_w2n_ro_icb_cmd_lock            ),
  .i0_icb_cmd_excl                (mst_g4_p0_w2n_ro_icb_cmd_excl            ),
  .i0_icb_cmd_xlen                (mst_g4_p0_w2n_ro_icb_cmd_xlen [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g4_p0_w2n_ro_icb_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (mst_g4_p0_w2n_ro_icb_cmd_modes [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g4_p0_w2n_ro_icb_cmd_dmode            ),
  .i0_icb_cmd_attri               (mst_g4_p0_w2n_ro_icb_cmd_attri [   2:   0]),
  .i0_icb_cmd_beat                (mst_g4_p0_w2n_ro_icb_cmd_beat [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g4_p0_w2n_ro_icb_cmd_usr  [   2:   0]),
  .i0_icb_rsp_ready               (mst_g4_p0_w2n_ro_icb_rsp_ready            ),
  .i0_icb_rsp_valid               (mst_g4_p0_w2n_ro_icb_rsp_valid            ),
  .i0_icb_rsp_err                 (mst_g4_p0_w2n_ro_icb_rsp_err             ),
  .i0_icb_rsp_excl_ok             (mst_g4_p0_w2n_ro_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g4_p0_w2n_ro_icb_rsp_rdata [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g4_p0_w2n_ro_icb_rsp_usr  [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_4_ro_icb_cmd_valid               ),
  .o_icb_cmd_ready                (mst_grp_4_ro_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (mst_grp_4_ro_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (mst_grp_4_ro_icb_cmd_read                ),
  .o_icb_cmd_addr                 (mst_grp_4_ro_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_4_ro_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_4_ro_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_4_ro_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_4_ro_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (mst_grp_4_ro_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (mst_grp_4_ro_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_4_ro_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_4_ro_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_4_ro_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (mst_grp_4_ro_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_4_ro_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_4_ro_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_4_ro_icb_rsp_ready               ),
  .o_icb_rsp_valid                (mst_grp_4_ro_icb_rsp_valid               ),
  .o_icb_rsp_err                  (mst_grp_4_ro_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (mst_grp_4_ro_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (mst_grp_4_ro_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_4_ro_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_mgrp4_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o4_wo_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g4_p0_w2n_wo_icb_cmd_valid            ),
  .i0_icb_cmd_ready               (mst_g4_p0_w2n_wo_icb_cmd_ready            ),
  .i0_icb_cmd_sel                 (mst_g4_p0_w2n_wo_icb_cmd_sel             ),
  .i0_icb_cmd_read                (mst_g4_p0_w2n_wo_icb_cmd_read            ),
  .i0_icb_cmd_addr                (mst_g4_p0_w2n_wo_icb_cmd_addr [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g4_p0_w2n_wo_icb_cmd_wdata [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g4_p0_w2n_wo_icb_cmd_wmask [   7:   0]),
  .i0_icb_cmd_size                (mst_g4_p0_w2n_wo_icb_cmd_size [   2:   0]),
  .i0_icb_cmd_lock                (mst_g4_p0_w2n_wo_icb_cmd_lock            ),
  .i0_icb_cmd_excl                (mst_g4_p0_w2n_wo_icb_cmd_excl            ),
  .i0_icb_cmd_xlen                (mst_g4_p0_w2n_wo_icb_cmd_xlen [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g4_p0_w2n_wo_icb_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (mst_g4_p0_w2n_wo_icb_cmd_modes [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g4_p0_w2n_wo_icb_cmd_dmode            ),
  .i0_icb_cmd_attri               (mst_g4_p0_w2n_wo_icb_cmd_attri [   2:   0]),
  .i0_icb_cmd_beat                (mst_g4_p0_w2n_wo_icb_cmd_beat [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g4_p0_w2n_wo_icb_cmd_usr  [   2:   0]),
  .i0_icb_rsp_ready               (mst_g4_p0_w2n_wo_icb_rsp_ready            ),
  .i0_icb_rsp_valid               (mst_g4_p0_w2n_wo_icb_rsp_valid            ),
  .i0_icb_rsp_err                 (mst_g4_p0_w2n_wo_icb_rsp_err             ),
  .i0_icb_rsp_excl_ok             (mst_g4_p0_w2n_wo_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g4_p0_w2n_wo_icb_rsp_rdata [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g4_p0_w2n_wo_icb_rsp_usr  [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_4_wo_icb_cmd_valid               ),
  .o_icb_cmd_ready                (mst_grp_4_wo_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (mst_grp_4_wo_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (mst_grp_4_wo_icb_cmd_read                ),
  .o_icb_cmd_addr                 (mst_grp_4_wo_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_4_wo_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_4_wo_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_4_wo_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_4_wo_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (mst_grp_4_wo_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (mst_grp_4_wo_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_4_wo_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_4_wo_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_4_wo_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (mst_grp_4_wo_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_4_wo_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_4_wo_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_4_wo_icb_rsp_ready               ),
  .o_icb_rsp_valid                (mst_grp_4_wo_icb_rsp_valid               ),
  .o_icb_rsp_err                  (mst_grp_4_wo_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (mst_grp_4_wo_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (mst_grp_4_wo_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_4_wo_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                mst_grp_5_icb_cmd_valid       ;
  wire                mst_grp_5_icb_cmd_ready       ;
  wire                mst_grp_5_icb_cmd_sel         ;
  wire                mst_grp_5_icb_cmd_read        ;
  wire    [  31:   0] mst_grp_5_icb_cmd_addr        ;
  wire    [  63:   0] mst_grp_5_icb_cmd_wdata       ;
  wire    [   7:   0] mst_grp_5_icb_cmd_wmask       ;
  wire    [   2:   0] mst_grp_5_icb_cmd_size        ;
  wire                mst_grp_5_icb_cmd_lock        ;
  wire                mst_grp_5_icb_cmd_excl        ;
  wire    [   7:   0] mst_grp_5_icb_cmd_xlen        ;
  wire    [   1:   0] mst_grp_5_icb_cmd_xburst      ;
  wire    [   1:   0] mst_grp_5_icb_cmd_modes       ;
  wire                mst_grp_5_icb_cmd_dmode       ;
  wire    [   2:   0] mst_grp_5_icb_cmd_attri       ;
  wire    [   1:   0] mst_grp_5_icb_cmd_beat        ;
  wire    [   2:   0] mst_grp_5_icb_cmd_usr         ;
  wire                mst_grp_5_icb_rsp_ready       ;
  wire                mst_grp_5_icb_rsp_valid       ;
  wire                mst_grp_5_icb_rsp_err         ;
  wire                mst_grp_5_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_grp_5_icb_rsp_rdata       ;
  wire    [   2:   0] mst_grp_5_icb_rsp_usr         ;
                 wire                mst_g5_p0_icb_cmd_valid       ;
  wire                mst_g5_p0_icb_cmd_ready       ;
  wire                mst_g5_p0_icb_cmd_sel         ;
  wire                mst_g5_p0_icb_cmd_read        ;
  wire    [  31:   0] mst_g5_p0_icb_cmd_addr        ;
  wire    [  63:   0] mst_g5_p0_icb_cmd_wdata       ;
  wire    [   7:   0] mst_g5_p0_icb_cmd_wmask       ;
  wire    [   2:   0] mst_g5_p0_icb_cmd_size        ;
  wire                mst_g5_p0_icb_cmd_lock        ;
  wire                mst_g5_p0_icb_cmd_excl        ;
  wire    [   7:   0] mst_g5_p0_icb_cmd_xlen        ;
  wire    [   1:   0] mst_g5_p0_icb_cmd_xburst      ;
  wire    [   1:   0] mst_g5_p0_icb_cmd_modes       ;
  wire                mst_g5_p0_icb_cmd_dmode       ;
  wire    [   2:   0] mst_g5_p0_icb_cmd_attri       ;
  wire    [   1:   0] mst_g5_p0_icb_cmd_beat        ;
  wire    [   2:   0] mst_g5_p0_icb_cmd_usr         ;
  wire                mst_g5_p0_icb_rsp_ready       ;
  wire                mst_g5_p0_icb_rsp_valid       ;
  wire                mst_g5_p0_icb_rsp_err         ;
  wire                mst_g5_p0_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_g5_p0_icb_rsp_rdata       ;
  wire    [   2:   0] mst_g5_p0_icb_rsp_usr         ;
                 wire                mst_g5_p0_w2n_icb_cmd_valid   ;
  wire                mst_g5_p0_w2n_icb_cmd_ready   ;
  wire                mst_g5_p0_w2n_icb_cmd_sel     ;
  wire                mst_g5_p0_w2n_icb_cmd_read    ;
  wire    [  31:   0] mst_g5_p0_w2n_icb_cmd_addr    ;
  wire    [  63:   0] mst_g5_p0_w2n_icb_cmd_wdata   ;
  wire    [   7:   0] mst_g5_p0_w2n_icb_cmd_wmask   ;
  wire    [   2:   0] mst_g5_p0_w2n_icb_cmd_size    ;
  wire                mst_g5_p0_w2n_icb_cmd_lock    ;
  wire                mst_g5_p0_w2n_icb_cmd_excl    ;
  wire    [   7:   0] mst_g5_p0_w2n_icb_cmd_xlen    ;
  wire    [   1:   0] mst_g5_p0_w2n_icb_cmd_xburst  ;
  wire    [   1:   0] mst_g5_p0_w2n_icb_cmd_modes   ;
  wire                mst_g5_p0_w2n_icb_cmd_dmode   ;
  wire    [   2:   0] mst_g5_p0_w2n_icb_cmd_attri   ;
  wire    [   1:   0] mst_g5_p0_w2n_icb_cmd_beat    ;
  wire    [   2:   0] mst_g5_p0_w2n_icb_cmd_usr     ;
  wire                mst_g5_p0_w2n_icb_rsp_ready   ;
  wire                mst_g5_p0_w2n_icb_rsp_valid   ;
  wire                mst_g5_p0_w2n_icb_rsp_err     ;
  wire                mst_g5_p0_w2n_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g5_p0_w2n_icb_rsp_rdata   ;
  wire    [   2:   0] mst_g5_p0_w2n_icb_rsp_usr     ;
    wire dummy_ahbl_bus_active;
               wire[3 -1:0] mst_g5_p0_icb_cmd_usr_pre;
               assign mst_g5_p0_icb_cmd_usr_pre = 3'b0;
               assign mst_g5_p0_icb_cmd_usr = mst_g5_p0_icb_cmd_usr_pre;
   e603_subsys_gnrl_usr_ahbl2ficb_ratio #(
       .SUPPORT_ICB_BURST(0),
      .SUPPORT_RATIO(0),
      .CMD_DP(2),
      .RSP_DP(2),
      .OUTS_CNT_W(7),
                .WR_EARLY_RETURN(1),
      .AW    (32),
      .DW    (64)  
    )u_dummy_ahbl_ahbl2ficb_ratio(
      .ratio_ahbl_clk_en(1'b1),
      .icb_clk_en   (1'b1),
      .ahbl2icb_ratio_active (dummy_ahbl_bus_active),
        .ahbl_htrans                    (dummy_ahbl_htrans             [   1:   0]),
  .ahbl_hwrite                    (dummy_ahbl_hwrite                        ),
  .ahbl_hmastlock                 (dummy_ahbl_hmastlock                     ),
  .ahbl_hsize                     (dummy_ahbl_hsize              [   2:   0]),
  .ahbl_hburst                    (dummy_ahbl_hburst             [   2:   0]),
  .ahbl_hprot                     (dummy_ahbl_hprot              [   3:   0]),
  .ahbl_hwdata                    (dummy_ahbl_hwdata             [  63:   0]),
  .ahbl_hrdata                    (dummy_ahbl_hrdata             [  63:   0]),
  .ahbl_hresp                     (dummy_ahbl_hresp              [   1:   0]),
  .ahbl_hready                    (dummy_ahbl_hready                        ),
      .ahbl_haddr(dummy_ahbl_haddr[32-1:0]),
      .ahbl_huser  (1'b0),
      .ahbl_hruser (),
       .icb_cmd_usr(),
       .icb_rsp_usr(1'b0),
        .icb_cmd_valid                  (mst_g5_p0_icb_cmd_valid                  ),
  .icb_cmd_ready                  (mst_g5_p0_icb_cmd_ready                  ),
  .icb_cmd_sel                    (mst_g5_p0_icb_cmd_sel                    ),
  .icb_cmd_read                   (mst_g5_p0_icb_cmd_read                   ),
  .icb_cmd_addr                   (mst_g5_p0_icb_cmd_addr        [  31:   0]),
  .icb_cmd_wdata                  (mst_g5_p0_icb_cmd_wdata       [  63:   0]),
  .icb_cmd_wmask                  (mst_g5_p0_icb_cmd_wmask       [   7:   0]),
  .icb_cmd_size                   (mst_g5_p0_icb_cmd_size        [   2:   0]),
  .icb_cmd_lock                   (mst_g5_p0_icb_cmd_lock                   ),
  .icb_cmd_excl                   (mst_g5_p0_icb_cmd_excl                   ),
  .icb_cmd_xlen                   (mst_g5_p0_icb_cmd_xlen        [   7:   0]),
  .icb_cmd_xburst                 (mst_g5_p0_icb_cmd_xburst      [   1:   0]),
  .icb_cmd_modes                  (mst_g5_p0_icb_cmd_modes       [   1:   0]),
  .icb_cmd_dmode                  (mst_g5_p0_icb_cmd_dmode                  ),
  .icb_cmd_attri                  (mst_g5_p0_icb_cmd_attri       [   2:   0]),
  .icb_cmd_beat                   (mst_g5_p0_icb_cmd_beat        [   1:   0]),
  .icb_rsp_ready                  (mst_g5_p0_icb_rsp_ready                  ),
  .icb_rsp_valid                  (mst_g5_p0_icb_rsp_valid                  ),
  .icb_rsp_err                    (mst_g5_p0_icb_rsp_err                    ),
  .icb_rsp_excl_ok                (mst_g5_p0_icb_rsp_excl_ok                ),
  .icb_rsp_rdata                  (mst_g5_p0_icb_rsp_rdata       [  63:   0]),
      .clk  (clk_fab),  
      .rst_n(rst_n)
    );
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g5_p0_icb_ficb_wconv(
        .i_icb_cmd_valid                (mst_g5_p0_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (mst_g5_p0_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (mst_g5_p0_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (mst_g5_p0_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (mst_g5_p0_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (mst_g5_p0_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (mst_g5_p0_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (mst_g5_p0_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (mst_g5_p0_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (mst_g5_p0_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (mst_g5_p0_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (mst_g5_p0_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (mst_g5_p0_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (mst_g5_p0_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (mst_g5_p0_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (mst_g5_p0_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (mst_g5_p0_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (mst_g5_p0_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (mst_g5_p0_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (mst_g5_p0_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (mst_g5_p0_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (mst_g5_p0_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (mst_g5_p0_icb_rsp_usr         [   2:   0]),
        .o_icb_cmd_valid                (mst_g5_p0_w2n_icb_cmd_valid              ),
  .o_icb_cmd_ready                (mst_g5_p0_w2n_icb_cmd_ready              ),
  .o_icb_cmd_sel                  (mst_g5_p0_w2n_icb_cmd_sel                ),
  .o_icb_cmd_read                 (mst_g5_p0_w2n_icb_cmd_read               ),
  .o_icb_cmd_addr                 (mst_g5_p0_w2n_icb_cmd_addr    [  31:   0]),
  .o_icb_cmd_wdata                (mst_g5_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .o_icb_cmd_wmask                (mst_g5_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .o_icb_cmd_size                 (mst_g5_p0_w2n_icb_cmd_size    [   2:   0]),
  .o_icb_cmd_lock                 (mst_g5_p0_w2n_icb_cmd_lock               ),
  .o_icb_cmd_excl                 (mst_g5_p0_w2n_icb_cmd_excl               ),
  .o_icb_cmd_xlen                 (mst_g5_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .o_icb_cmd_xburst               (mst_g5_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .o_icb_cmd_modes                (mst_g5_p0_w2n_icb_cmd_modes   [   1:   0]),
  .o_icb_cmd_dmode                (mst_g5_p0_w2n_icb_cmd_dmode              ),
  .o_icb_cmd_attri                (mst_g5_p0_w2n_icb_cmd_attri   [   2:   0]),
  .o_icb_cmd_beat                 (mst_g5_p0_w2n_icb_cmd_beat    [   1:   0]),
  .o_icb_cmd_usr                  (mst_g5_p0_w2n_icb_cmd_usr     [   2:   0]),
  .o_icb_rsp_ready                (mst_g5_p0_w2n_icb_rsp_ready              ),
  .o_icb_rsp_valid                (mst_g5_p0_w2n_icb_rsp_valid              ),
  .o_icb_rsp_err                  (mst_g5_p0_w2n_icb_rsp_err                ),
  .o_icb_rsp_excl_ok              (mst_g5_p0_w2n_icb_rsp_excl_ok            ),
  .o_icb_rsp_rdata                (mst_g5_p0_w2n_icb_rsp_rdata   [  63:   0]),
  .o_icb_rsp_usr                  (mst_g5_p0_w2n_icb_rsp_usr     [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   e603_subsys_mgrp5_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o5_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g5_p0_w2n_icb_cmd_valid              ),
  .i0_icb_cmd_ready               (mst_g5_p0_w2n_icb_cmd_ready              ),
  .i0_icb_cmd_sel                 (mst_g5_p0_w2n_icb_cmd_sel                ),
  .i0_icb_cmd_read                (mst_g5_p0_w2n_icb_cmd_read               ),
  .i0_icb_cmd_addr                (mst_g5_p0_w2n_icb_cmd_addr    [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g5_p0_w2n_icb_cmd_wdata   [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g5_p0_w2n_icb_cmd_wmask   [   7:   0]),
  .i0_icb_cmd_size                (mst_g5_p0_w2n_icb_cmd_size    [   2:   0]),
  .i0_icb_cmd_lock                (mst_g5_p0_w2n_icb_cmd_lock               ),
  .i0_icb_cmd_excl                (mst_g5_p0_w2n_icb_cmd_excl               ),
  .i0_icb_cmd_xlen                (mst_g5_p0_w2n_icb_cmd_xlen    [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g5_p0_w2n_icb_cmd_xburst  [   1:   0]),
  .i0_icb_cmd_modes               (mst_g5_p0_w2n_icb_cmd_modes   [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g5_p0_w2n_icb_cmd_dmode              ),
  .i0_icb_cmd_attri               (mst_g5_p0_w2n_icb_cmd_attri   [   2:   0]),
  .i0_icb_cmd_beat                (mst_g5_p0_w2n_icb_cmd_beat    [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g5_p0_w2n_icb_cmd_usr     [   2:   0]),
  .i0_icb_rsp_ready               (mst_g5_p0_w2n_icb_rsp_ready              ),
  .i0_icb_rsp_valid               (mst_g5_p0_w2n_icb_rsp_valid              ),
  .i0_icb_rsp_err                 (mst_g5_p0_w2n_icb_rsp_err                ),
  .i0_icb_rsp_excl_ok             (mst_g5_p0_w2n_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g5_p0_w2n_icb_rsp_rdata   [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g5_p0_w2n_icb_rsp_usr     [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_5_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (mst_grp_5_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (mst_grp_5_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (mst_grp_5_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (mst_grp_5_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_5_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_5_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_5_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_5_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (mst_grp_5_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (mst_grp_5_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_5_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_5_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_5_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (mst_grp_5_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_5_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_5_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_5_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (mst_grp_5_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (mst_grp_5_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (mst_grp_5_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (mst_grp_5_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_5_icb_rsp_usr         [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                mst_grp_6_ro_icb_cmd_valid    ;
  wire                mst_grp_6_ro_icb_cmd_ready    ;
  wire                mst_grp_6_ro_icb_cmd_sel      ;
  wire                mst_grp_6_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_6_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_6_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_6_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_6_ro_icb_cmd_size     ;
  wire                mst_grp_6_ro_icb_cmd_lock     ;
  wire                mst_grp_6_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_6_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_6_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_6_ro_icb_cmd_modes    ;
  wire                mst_grp_6_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_6_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_6_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_6_ro_icb_cmd_usr      ;
  wire                mst_grp_6_ro_icb_rsp_ready    ;
  wire                mst_grp_6_ro_icb_rsp_valid    ;
  wire                mst_grp_6_ro_icb_rsp_err      ;
  wire                mst_grp_6_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_6_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_6_ro_icb_rsp_usr      ;
      wire                mst_grp_6_wo_icb_cmd_valid    ;
  wire                mst_grp_6_wo_icb_cmd_ready    ;
  wire                mst_grp_6_wo_icb_cmd_sel      ;
  wire                mst_grp_6_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_6_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_6_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_6_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_6_wo_icb_cmd_size     ;
  wire                mst_grp_6_wo_icb_cmd_lock     ;
  wire                mst_grp_6_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_6_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_6_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_6_wo_icb_cmd_modes    ;
  wire                mst_grp_6_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_6_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_6_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_6_wo_icb_cmd_usr      ;
  wire                mst_grp_6_wo_icb_rsp_ready    ;
  wire                mst_grp_6_wo_icb_rsp_valid    ;
  wire                mst_grp_6_wo_icb_rsp_err      ;
  wire                mst_grp_6_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_6_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_6_wo_icb_rsp_usr      ;
                 wire                mst_g6_p0_icb_cmd_valid       ;
  wire                mst_g6_p0_icb_cmd_ready       ;
  wire                mst_g6_p0_icb_cmd_sel         ;
  wire                mst_g6_p0_icb_cmd_read        ;
  wire    [  31:   0] mst_g6_p0_icb_cmd_addr        ;
  wire    [  63:   0] mst_g6_p0_icb_cmd_wdata       ;
  wire    [   7:   0] mst_g6_p0_icb_cmd_wmask       ;
  wire    [   2:   0] mst_g6_p0_icb_cmd_size        ;
  wire                mst_g6_p0_icb_cmd_lock        ;
  wire                mst_g6_p0_icb_cmd_excl        ;
  wire    [   7:   0] mst_g6_p0_icb_cmd_xlen        ;
  wire    [   1:   0] mst_g6_p0_icb_cmd_xburst      ;
  wire    [   1:   0] mst_g6_p0_icb_cmd_modes       ;
  wire                mst_g6_p0_icb_cmd_dmode       ;
  wire    [   2:   0] mst_g6_p0_icb_cmd_attri       ;
  wire    [   1:   0] mst_g6_p0_icb_cmd_beat        ;
  wire    [   2:   0] mst_g6_p0_icb_cmd_usr         ;
  wire                mst_g6_p0_icb_rsp_ready       ;
  wire                mst_g6_p0_icb_rsp_valid       ;
  wire                mst_g6_p0_icb_rsp_err         ;
  wire                mst_g6_p0_icb_rsp_excl_ok     ;
  wire    [  63:   0] mst_g6_p0_icb_rsp_rdata       ;
  wire    [   2:   0] mst_g6_p0_icb_rsp_usr         ;
                 wire                mst_g6_p0_w2n_ro_icb_cmd_valid ;
  wire                mst_g6_p0_w2n_ro_icb_cmd_ready ;
  wire                mst_g6_p0_w2n_ro_icb_cmd_sel  ;
  wire                mst_g6_p0_w2n_ro_icb_cmd_read ;
  wire    [  31:   0] mst_g6_p0_w2n_ro_icb_cmd_addr ;
  wire    [  63:   0] mst_g6_p0_w2n_ro_icb_cmd_wdata ;
  wire    [   7:   0] mst_g6_p0_w2n_ro_icb_cmd_wmask ;
  wire    [   2:   0] mst_g6_p0_w2n_ro_icb_cmd_size ;
  wire                mst_g6_p0_w2n_ro_icb_cmd_lock ;
  wire                mst_g6_p0_w2n_ro_icb_cmd_excl ;
  wire    [   7:   0] mst_g6_p0_w2n_ro_icb_cmd_xlen ;
  wire    [   1:   0] mst_g6_p0_w2n_ro_icb_cmd_xburst ;
  wire    [   1:   0] mst_g6_p0_w2n_ro_icb_cmd_modes ;
  wire                mst_g6_p0_w2n_ro_icb_cmd_dmode ;
  wire    [   2:   0] mst_g6_p0_w2n_ro_icb_cmd_attri ;
  wire    [   1:   0] mst_g6_p0_w2n_ro_icb_cmd_beat ;
  wire    [   2:   0] mst_g6_p0_w2n_ro_icb_cmd_usr  ;
  wire                mst_g6_p0_w2n_ro_icb_rsp_ready ;
  wire                mst_g6_p0_w2n_ro_icb_rsp_valid ;
  wire                mst_g6_p0_w2n_ro_icb_rsp_err  ;
  wire                mst_g6_p0_w2n_ro_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g6_p0_w2n_ro_icb_rsp_rdata ;
  wire    [   2:   0] mst_g6_p0_w2n_ro_icb_rsp_usr  ;
                 wire                mst_g6_p0_w2n_wo_icb_cmd_valid ;
  wire                mst_g6_p0_w2n_wo_icb_cmd_ready ;
  wire                mst_g6_p0_w2n_wo_icb_cmd_sel  ;
  wire                mst_g6_p0_w2n_wo_icb_cmd_read ;
  wire    [  31:   0] mst_g6_p0_w2n_wo_icb_cmd_addr ;
  wire    [  63:   0] mst_g6_p0_w2n_wo_icb_cmd_wdata ;
  wire    [   7:   0] mst_g6_p0_w2n_wo_icb_cmd_wmask ;
  wire    [   2:   0] mst_g6_p0_w2n_wo_icb_cmd_size ;
  wire                mst_g6_p0_w2n_wo_icb_cmd_lock ;
  wire                mst_g6_p0_w2n_wo_icb_cmd_excl ;
  wire    [   7:   0] mst_g6_p0_w2n_wo_icb_cmd_xlen ;
  wire    [   1:   0] mst_g6_p0_w2n_wo_icb_cmd_xburst ;
  wire    [   1:   0] mst_g6_p0_w2n_wo_icb_cmd_modes ;
  wire                mst_g6_p0_w2n_wo_icb_cmd_dmode ;
  wire    [   2:   0] mst_g6_p0_w2n_wo_icb_cmd_attri ;
  wire    [   1:   0] mst_g6_p0_w2n_wo_icb_cmd_beat ;
  wire    [   2:   0] mst_g6_p0_w2n_wo_icb_cmd_usr  ;
  wire                mst_g6_p0_w2n_wo_icb_rsp_ready ;
  wire                mst_g6_p0_w2n_wo_icb_rsp_valid ;
  wire                mst_g6_p0_w2n_wo_icb_rsp_err  ;
  wire                mst_g6_p0_w2n_wo_icb_rsp_excl_ok ;
  wire    [  63:   0] mst_g6_p0_w2n_wo_icb_rsp_rdata ;
  wire    [   2:   0] mst_g6_p0_w2n_wo_icb_rsp_usr  ;
    wire eth_axi_bus_active;
                 wire                mst_g6_p0_ro_icb_cmd_valid    ;
  wire                mst_g6_p0_ro_icb_cmd_ready    ;
  wire                mst_g6_p0_ro_icb_cmd_sel      ;
  wire                mst_g6_p0_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_g6_p0_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_g6_p0_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_g6_p0_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_g6_p0_ro_icb_cmd_size     ;
  wire                mst_g6_p0_ro_icb_cmd_lock     ;
  wire                mst_g6_p0_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_g6_p0_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_g6_p0_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_g6_p0_ro_icb_cmd_modes    ;
  wire                mst_g6_p0_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_g6_p0_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_g6_p0_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_g6_p0_ro_icb_cmd_usr      ;
  wire                mst_g6_p0_ro_icb_rsp_ready    ;
  wire                mst_g6_p0_ro_icb_rsp_valid    ;
  wire                mst_g6_p0_ro_icb_rsp_err      ;
  wire                mst_g6_p0_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_g6_p0_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_g6_p0_ro_icb_rsp_usr      ;
    wire mst_g6_p0_ro_icb_bus_active;
                              wire[3-1:0] mst_g6_p0_ro_icb_cmd_usr_pre;
               assign mst_g6_p0_ro_icb_cmd_usr = mst_g6_p0_ro_icb_cmd_usr_pre;
  e603_subsys_gnrl_axi2ficb_read_async # (
      .ID_W(1),
    .SYNC_DP       (2),
    .ASYNC_FIFO    (1),
    .ASYNC_FIFO_DP (8),
    .ASYNC_FIFO_DP_PTR_W (3),
      .AW(32),
      .DW(64), 
      .MW(64/8), 
      .FIFO_OUTS_NUM (64),
      .USR_W (3)
    )u_eth_axi_axi2ficb_read(
  .reset_flag_r  (1'b0),
      .axi_arvalid                    (eth_axi_arvalid                          ),
  .axi_arready                    (eth_axi_arready                          ),
  .axi_arlen                      (eth_axi_arlen                 [   7:   0]),
  .axi_arsize                     (eth_axi_arsize                [   2:   0]),
  .axi_arburst                    (eth_axi_arburst               [   1:   0]),
  .axi_arlock                     (eth_axi_arlock                           ),
  .axi_arcache                    (eth_axi_arcache               [   3:   0]),
  .axi_arprot                     (eth_axi_arprot                [   2:   0]),
  .axi_rready                     (eth_axi_rready                           ),
  .axi_rvalid                     (eth_axi_rvalid                           ),
  .axi_rdata                      (eth_axi_rdata                 [  63:   0]),
  .axi_rresp                      (eth_axi_rresp                 [   1:   0]),
  .axi_rlast                      (eth_axi_rlast                            ),
      .axi_araddr(eth_axi_araddr[32-1:0]),
      .axi_aruser(3'b0),
      .axi_ruser(),
      .axi_arid(1'b0),
      .axi_rid (),
        .icb_rcmd_valid                 (mst_g6_p0_ro_icb_cmd_valid               ),
  .icb_rcmd_ready                 (mst_g6_p0_ro_icb_cmd_ready               ),
  .icb_rcmd_sel                   (mst_g6_p0_ro_icb_cmd_sel                 ),
  .icb_rcmd_read                  (mst_g6_p0_ro_icb_cmd_read                ),
  .icb_rcmd_addr                  (mst_g6_p0_ro_icb_cmd_addr     [  31:   0]),
  .icb_rcmd_wdata                 (mst_g6_p0_ro_icb_cmd_wdata    [  63:   0]),
  .icb_rcmd_wmask                 (mst_g6_p0_ro_icb_cmd_wmask    [   7:   0]),
  .icb_rcmd_size                  (mst_g6_p0_ro_icb_cmd_size     [   2:   0]),
  .icb_rcmd_excl                  (mst_g6_p0_ro_icb_cmd_excl                ),
  .icb_rcmd_xlen                  (mst_g6_p0_ro_icb_cmd_xlen     [   7:   0]),
  .icb_rcmd_xburst                (mst_g6_p0_ro_icb_cmd_xburst   [   1:   0]),
  .icb_rcmd_modes                 (mst_g6_p0_ro_icb_cmd_modes    [   1:   0]),
  .icb_rcmd_dmode                 (mst_g6_p0_ro_icb_cmd_dmode               ),
  .icb_rcmd_attri                 (mst_g6_p0_ro_icb_cmd_attri    [   2:   0]),
  .icb_rcmd_beat                  (mst_g6_p0_ro_icb_cmd_beat     [   1:   0]),
  .icb_rrsp_ready                 (mst_g6_p0_ro_icb_rsp_ready               ),
  .icb_rrsp_valid                 (mst_g6_p0_ro_icb_rsp_valid               ),
  .icb_rrsp_err                   (mst_g6_p0_ro_icb_rsp_err                 ),
  .icb_rrsp_excl_ok               (mst_g6_p0_ro_icb_rsp_excl_ok             ),
  .icb_rrsp_rdata                 (mst_g6_p0_ro_icb_rsp_rdata    [  63:   0]),
      .icb_rcmd_usr(mst_g6_p0_ro_icb_cmd_usr_pre),
      .icb_rrsp_usr(mst_g6_p0_ro_icb_rsp_usr[3-1:0]),
      .axi2icb_read_axi_active (),
      .axi2icb_read_icb_active (mst_g6_p0_ro_icb_bus_active),
      .async_axi_clk  (eth_axi_clk  ),
      .async_axi_rst_n(eth_axi_rst_n_sync_4port), 
      .icb_clk  (clk),
      .icb_rst_n(eth_axi_rst_n_sync_4fab)
    );
    assign mst_g6_p0_ro_icb_cmd_lock = 1'b0;
                 wire                mst_g6_p0_wo_icb_cmd_valid    ;
  wire                mst_g6_p0_wo_icb_cmd_ready    ;
  wire                mst_g6_p0_wo_icb_cmd_sel      ;
  wire                mst_g6_p0_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_g6_p0_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_g6_p0_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_g6_p0_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_g6_p0_wo_icb_cmd_size     ;
  wire                mst_g6_p0_wo_icb_cmd_lock     ;
  wire                mst_g6_p0_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_g6_p0_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_g6_p0_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_g6_p0_wo_icb_cmd_modes    ;
  wire                mst_g6_p0_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_g6_p0_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_g6_p0_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_g6_p0_wo_icb_cmd_usr      ;
  wire                mst_g6_p0_wo_icb_rsp_ready    ;
  wire                mst_g6_p0_wo_icb_rsp_valid    ;
  wire                mst_g6_p0_wo_icb_rsp_err      ;
  wire                mst_g6_p0_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_g6_p0_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_g6_p0_wo_icb_rsp_usr      ;
    wire mst_g6_p0_wo_icb_bus_active;
                              wire[3-1:0] mst_g6_p0_wo_icb_cmd_usr_pre;
               assign mst_g6_p0_wo_icb_cmd_usr = mst_g6_p0_wo_icb_cmd_usr_pre;
  e603_subsys_gnrl_axi2ficb_write_async # (
      .ID_W(1),
    .SYNC_DP       (2),
    .ASYNC_FIFO    (1),
    .ASYNC_FIFO_DP (8),
    .ASYNC_FIFO_DP_PTR_W (3),
      .AW(32),
      .DW(64), 
      .MW(64/8), 
      .FIFO_OUTS_NUM (64),
      .USR_W (3)
    )u_mst_g6_p0_wo_icb_axi2ficb_write(
  .reset_flag_r  (1'b0),
      .axi_awvalid                    (eth_axi_awvalid                          ),
  .axi_awready                    (eth_axi_awready                          ),
  .axi_awlen                      (eth_axi_awlen                 [   7:   0]),
  .axi_awsize                     (eth_axi_awsize                [   2:   0]),
  .axi_awburst                    (eth_axi_awburst               [   1:   0]),
  .axi_awlock                     (eth_axi_awlock                           ),
  .axi_awcache                    (eth_axi_awcache               [   3:   0]),
  .axi_awprot                     (eth_axi_awprot                [   2:   0]),
  .axi_bready                     (eth_axi_bready                           ),
  .axi_bvalid                     (eth_axi_bvalid                           ),
  .axi_bresp                      (eth_axi_bresp                 [   1:   0]),
  .axi_wready                     (eth_axi_wready                           ),
  .axi_wvalid                     (eth_axi_wvalid                           ),
  .axi_wdata                      (eth_axi_wdata                 [  63:   0]),
  .axi_wstrb                      (eth_axi_wstrb                 [   7:   0]),
  .axi_wlast                      (eth_axi_wlast                            ),
      .axi_awaddr(eth_axi_awaddr[32-1:0]),
      .axi_awuser(3'b0),
      .axi_buser(),
      .axi_awid(1'b0),
      .axi_bid (),
        .icb_wcmd_valid                 (mst_g6_p0_wo_icb_cmd_valid               ),
  .icb_wcmd_ready                 (mst_g6_p0_wo_icb_cmd_ready               ),
  .icb_wcmd_sel                   (mst_g6_p0_wo_icb_cmd_sel                 ),
  .icb_wcmd_read                  (mst_g6_p0_wo_icb_cmd_read                ),
  .icb_wcmd_addr                  (mst_g6_p0_wo_icb_cmd_addr     [  31:   0]),
  .icb_wcmd_wdata                 (mst_g6_p0_wo_icb_cmd_wdata    [  63:   0]),
  .icb_wcmd_wmask                 (mst_g6_p0_wo_icb_cmd_wmask    [   7:   0]),
  .icb_wcmd_size                  (mst_g6_p0_wo_icb_cmd_size     [   2:   0]),
  .icb_wcmd_lock                  (mst_g6_p0_wo_icb_cmd_lock                ),
  .icb_wcmd_excl                  (mst_g6_p0_wo_icb_cmd_excl                ),
  .icb_wcmd_xlen                  (mst_g6_p0_wo_icb_cmd_xlen     [   7:   0]),
  .icb_wcmd_xburst                (mst_g6_p0_wo_icb_cmd_xburst   [   1:   0]),
  .icb_wcmd_modes                 (mst_g6_p0_wo_icb_cmd_modes    [   1:   0]),
  .icb_wcmd_dmode                 (mst_g6_p0_wo_icb_cmd_dmode               ),
  .icb_wcmd_attri                 (mst_g6_p0_wo_icb_cmd_attri    [   2:   0]),
  .icb_wcmd_beat                  (mst_g6_p0_wo_icb_cmd_beat     [   1:   0]),
  .icb_wrsp_ready                 (mst_g6_p0_wo_icb_rsp_ready               ),
  .icb_wrsp_valid                 (mst_g6_p0_wo_icb_rsp_valid               ),
  .icb_wrsp_err                   (mst_g6_p0_wo_icb_rsp_err                 ),
  .icb_wrsp_excl_ok               (mst_g6_p0_wo_icb_rsp_excl_ok             ),
      .icb_wcmd_usr(mst_g6_p0_wo_icb_cmd_usr_pre),
      .icb_wrsp_usr(mst_g6_p0_wo_icb_rsp_usr[3-1:0]),
      .axi2icb_write_axi_active (),
      .axi2icb_write_icb_active (mst_g6_p0_wo_icb_bus_active),
      .async_axi_clk  (eth_axi_clk  ),
      .async_axi_rst_n(eth_axi_rst_n_sync_4port), 
      .icb_clk  (clk),
      .icb_rst_n(eth_axi_rst_n_sync_4fab)
    );
   assign eth_axi_bus_active = 1'b0
                     | mst_g6_p0_ro_icb_bus_active
                     | mst_g6_p0_wo_icb_bus_active
                 ;
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g6_p0_ro_icb_ficb_wconv(
      .i_icb_cmd_read(1'b1),
                .i_icb_cmd_wdata (64'b0),
                .i_icb_cmd_wmask (8'b0),
        .i_icb_cmd_valid                (mst_g6_p0_ro_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_g6_p0_ro_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_g6_p0_ro_icb_cmd_sel                 ),
  .i_icb_cmd_addr                 (mst_g6_p0_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_size                 (mst_g6_p0_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_g6_p0_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_g6_p0_ro_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_g6_p0_ro_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_g6_p0_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_g6_p0_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_g6_p0_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_g6_p0_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_g6_p0_ro_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_g6_p0_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_g6_p0_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_g6_p0_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_g6_p0_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_g6_p0_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_g6_p0_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_g6_p0_ro_icb_rsp_usr      [   2:   0]),
        .o_icb_cmd_valid                (mst_g6_p0_w2n_ro_icb_cmd_valid            ),
  .o_icb_cmd_ready                (mst_g6_p0_w2n_ro_icb_cmd_ready            ),
  .o_icb_cmd_sel                  (mst_g6_p0_w2n_ro_icb_cmd_sel             ),
  .o_icb_cmd_read                 (mst_g6_p0_w2n_ro_icb_cmd_read            ),
  .o_icb_cmd_addr                 (mst_g6_p0_w2n_ro_icb_cmd_addr [  31:   0]),
  .o_icb_cmd_wdata                (mst_g6_p0_w2n_ro_icb_cmd_wdata [  63:   0]),
  .o_icb_cmd_wmask                (mst_g6_p0_w2n_ro_icb_cmd_wmask [   7:   0]),
  .o_icb_cmd_size                 (mst_g6_p0_w2n_ro_icb_cmd_size [   2:   0]),
  .o_icb_cmd_lock                 (mst_g6_p0_w2n_ro_icb_cmd_lock            ),
  .o_icb_cmd_excl                 (mst_g6_p0_w2n_ro_icb_cmd_excl            ),
  .o_icb_cmd_xlen                 (mst_g6_p0_w2n_ro_icb_cmd_xlen [   7:   0]),
  .o_icb_cmd_xburst               (mst_g6_p0_w2n_ro_icb_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (mst_g6_p0_w2n_ro_icb_cmd_modes [   1:   0]),
  .o_icb_cmd_dmode                (mst_g6_p0_w2n_ro_icb_cmd_dmode            ),
  .o_icb_cmd_attri                (mst_g6_p0_w2n_ro_icb_cmd_attri [   2:   0]),
  .o_icb_cmd_beat                 (mst_g6_p0_w2n_ro_icb_cmd_beat [   1:   0]),
  .o_icb_cmd_usr                  (mst_g6_p0_w2n_ro_icb_cmd_usr  [   2:   0]),
  .o_icb_rsp_ready                (mst_g6_p0_w2n_ro_icb_rsp_ready            ),
  .o_icb_rsp_valid                (mst_g6_p0_w2n_ro_icb_rsp_valid            ),
  .o_icb_rsp_err                  (mst_g6_p0_w2n_ro_icb_rsp_err             ),
  .o_icb_rsp_excl_ok              (mst_g6_p0_w2n_ro_icb_rsp_excl_ok            ),
  .o_icb_rsp_rdata                (mst_g6_p0_w2n_ro_icb_rsp_rdata [  63:   0]),
  .o_icb_rsp_usr                  (mst_g6_p0_w2n_ro_icb_rsp_usr  [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .RSP_CHECK_CMD_OUTS(RSP_CHECK_CMD_OUTS),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .AW    (32),
      .ZEROCYC_RSP   (0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .FIFO_OUTS_NUM (64),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_mst_g6_p0_wo_icb_ficb_wconv(
        .i_icb_cmd_valid                (mst_g6_p0_wo_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_g6_p0_wo_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_g6_p0_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_g6_p0_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_g6_p0_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_g6_p0_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_g6_p0_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_g6_p0_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_g6_p0_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_g6_p0_wo_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_g6_p0_wo_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_g6_p0_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_g6_p0_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_g6_p0_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_g6_p0_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_g6_p0_wo_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_g6_p0_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_g6_p0_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_g6_p0_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_g6_p0_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_g6_p0_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_g6_p0_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_g6_p0_wo_icb_rsp_usr      [   2:   0]),
                .o_icb_rsp_rdata (64'b0),
        .o_icb_cmd_valid                (mst_g6_p0_w2n_wo_icb_cmd_valid            ),
  .o_icb_cmd_ready                (mst_g6_p0_w2n_wo_icb_cmd_ready            ),
  .o_icb_cmd_sel                  (mst_g6_p0_w2n_wo_icb_cmd_sel             ),
  .o_icb_cmd_read                 (mst_g6_p0_w2n_wo_icb_cmd_read            ),
  .o_icb_cmd_addr                 (mst_g6_p0_w2n_wo_icb_cmd_addr [  31:   0]),
  .o_icb_cmd_wdata                (mst_g6_p0_w2n_wo_icb_cmd_wdata [  63:   0]),
  .o_icb_cmd_wmask                (mst_g6_p0_w2n_wo_icb_cmd_wmask [   7:   0]),
  .o_icb_cmd_size                 (mst_g6_p0_w2n_wo_icb_cmd_size [   2:   0]),
  .o_icb_cmd_lock                 (mst_g6_p0_w2n_wo_icb_cmd_lock            ),
  .o_icb_cmd_excl                 (mst_g6_p0_w2n_wo_icb_cmd_excl            ),
  .o_icb_cmd_xlen                 (mst_g6_p0_w2n_wo_icb_cmd_xlen [   7:   0]),
  .o_icb_cmd_xburst               (mst_g6_p0_w2n_wo_icb_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (mst_g6_p0_w2n_wo_icb_cmd_modes [   1:   0]),
  .o_icb_cmd_dmode                (mst_g6_p0_w2n_wo_icb_cmd_dmode            ),
  .o_icb_cmd_attri                (mst_g6_p0_w2n_wo_icb_cmd_attri [   2:   0]),
  .o_icb_cmd_beat                 (mst_g6_p0_w2n_wo_icb_cmd_beat [   1:   0]),
  .o_icb_cmd_usr                  (mst_g6_p0_w2n_wo_icb_cmd_usr  [   2:   0]),
  .o_icb_rsp_ready                (mst_g6_p0_w2n_wo_icb_rsp_ready            ),
  .o_icb_rsp_valid                (mst_g6_p0_w2n_wo_icb_rsp_valid            ),
  .o_icb_rsp_err                  (mst_g6_p0_w2n_wo_icb_rsp_err             ),
  .o_icb_rsp_excl_ok              (mst_g6_p0_w2n_wo_icb_rsp_excl_ok            ),
  .o_icb_rsp_usr                  (mst_g6_p0_w2n_wo_icb_rsp_usr  [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
   e603_subsys_mgrp6_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o6_ro_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g6_p0_w2n_ro_icb_cmd_valid            ),
  .i0_icb_cmd_ready               (mst_g6_p0_w2n_ro_icb_cmd_ready            ),
  .i0_icb_cmd_sel                 (mst_g6_p0_w2n_ro_icb_cmd_sel             ),
  .i0_icb_cmd_read                (mst_g6_p0_w2n_ro_icb_cmd_read            ),
  .i0_icb_cmd_addr                (mst_g6_p0_w2n_ro_icb_cmd_addr [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g6_p0_w2n_ro_icb_cmd_wdata [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g6_p0_w2n_ro_icb_cmd_wmask [   7:   0]),
  .i0_icb_cmd_size                (mst_g6_p0_w2n_ro_icb_cmd_size [   2:   0]),
  .i0_icb_cmd_lock                (mst_g6_p0_w2n_ro_icb_cmd_lock            ),
  .i0_icb_cmd_excl                (mst_g6_p0_w2n_ro_icb_cmd_excl            ),
  .i0_icb_cmd_xlen                (mst_g6_p0_w2n_ro_icb_cmd_xlen [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g6_p0_w2n_ro_icb_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (mst_g6_p0_w2n_ro_icb_cmd_modes [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g6_p0_w2n_ro_icb_cmd_dmode            ),
  .i0_icb_cmd_attri               (mst_g6_p0_w2n_ro_icb_cmd_attri [   2:   0]),
  .i0_icb_cmd_beat                (mst_g6_p0_w2n_ro_icb_cmd_beat [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g6_p0_w2n_ro_icb_cmd_usr  [   2:   0]),
  .i0_icb_rsp_ready               (mst_g6_p0_w2n_ro_icb_rsp_ready            ),
  .i0_icb_rsp_valid               (mst_g6_p0_w2n_ro_icb_rsp_valid            ),
  .i0_icb_rsp_err                 (mst_g6_p0_w2n_ro_icb_rsp_err             ),
  .i0_icb_rsp_excl_ok             (mst_g6_p0_w2n_ro_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g6_p0_w2n_ro_icb_rsp_rdata [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g6_p0_w2n_ro_icb_rsp_usr  [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_6_ro_icb_cmd_valid               ),
  .o_icb_cmd_ready                (mst_grp_6_ro_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (mst_grp_6_ro_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (mst_grp_6_ro_icb_cmd_read                ),
  .o_icb_cmd_addr                 (mst_grp_6_ro_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_6_ro_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_6_ro_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_6_ro_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_6_ro_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (mst_grp_6_ro_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (mst_grp_6_ro_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_6_ro_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_6_ro_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_6_ro_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (mst_grp_6_ro_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_6_ro_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_6_ro_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_6_ro_icb_rsp_ready               ),
  .o_icb_rsp_valid                (mst_grp_6_ro_icb_rsp_valid               ),
  .o_icb_rsp_err                  (mst_grp_6_ro_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (mst_grp_6_ro_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (mst_grp_6_ro_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_6_ro_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_mgrp6_ficbnto1_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .SUPPORT_LOCK(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ARBT_SCHEME            (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP   (0),
      .ARBT_FIFO_OUTS_NUM  (64  ),
      .ARBT_FIFO_OUTS_CNT_W(7),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_arbt_o6_wo_icb(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (),
                    .i0_icb_cmd_valid               (mst_g6_p0_w2n_wo_icb_cmd_valid            ),
  .i0_icb_cmd_ready               (mst_g6_p0_w2n_wo_icb_cmd_ready            ),
  .i0_icb_cmd_sel                 (mst_g6_p0_w2n_wo_icb_cmd_sel             ),
  .i0_icb_cmd_read                (mst_g6_p0_w2n_wo_icb_cmd_read            ),
  .i0_icb_cmd_addr                (mst_g6_p0_w2n_wo_icb_cmd_addr [  31:   0]),
  .i0_icb_cmd_wdata               (mst_g6_p0_w2n_wo_icb_cmd_wdata [  63:   0]),
  .i0_icb_cmd_wmask               (mst_g6_p0_w2n_wo_icb_cmd_wmask [   7:   0]),
  .i0_icb_cmd_size                (mst_g6_p0_w2n_wo_icb_cmd_size [   2:   0]),
  .i0_icb_cmd_lock                (mst_g6_p0_w2n_wo_icb_cmd_lock            ),
  .i0_icb_cmd_excl                (mst_g6_p0_w2n_wo_icb_cmd_excl            ),
  .i0_icb_cmd_xlen                (mst_g6_p0_w2n_wo_icb_cmd_xlen [   7:   0]),
  .i0_icb_cmd_xburst              (mst_g6_p0_w2n_wo_icb_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (mst_g6_p0_w2n_wo_icb_cmd_modes [   1:   0]),
  .i0_icb_cmd_dmode               (mst_g6_p0_w2n_wo_icb_cmd_dmode            ),
  .i0_icb_cmd_attri               (mst_g6_p0_w2n_wo_icb_cmd_attri [   2:   0]),
  .i0_icb_cmd_beat                (mst_g6_p0_w2n_wo_icb_cmd_beat [   1:   0]),
  .i0_icb_cmd_usr                 (mst_g6_p0_w2n_wo_icb_cmd_usr  [   2:   0]),
  .i0_icb_rsp_ready               (mst_g6_p0_w2n_wo_icb_rsp_ready            ),
  .i0_icb_rsp_valid               (mst_g6_p0_w2n_wo_icb_rsp_valid            ),
  .i0_icb_rsp_err                 (mst_g6_p0_w2n_wo_icb_rsp_err             ),
  .i0_icb_rsp_excl_ok             (mst_g6_p0_w2n_wo_icb_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (mst_g6_p0_w2n_wo_icb_rsp_rdata [  63:   0]),
  .i0_icb_rsp_usr                 (mst_g6_p0_w2n_wo_icb_rsp_usr  [   2:   0]),
      .o_icb_cmd_valid                (mst_grp_6_wo_icb_cmd_valid               ),
  .o_icb_cmd_ready                (mst_grp_6_wo_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (mst_grp_6_wo_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (mst_grp_6_wo_icb_cmd_read                ),
  .o_icb_cmd_addr                 (mst_grp_6_wo_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (mst_grp_6_wo_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (mst_grp_6_wo_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (mst_grp_6_wo_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (mst_grp_6_wo_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (mst_grp_6_wo_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (mst_grp_6_wo_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (mst_grp_6_wo_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (mst_grp_6_wo_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (mst_grp_6_wo_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (mst_grp_6_wo_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (mst_grp_6_wo_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (mst_grp_6_wo_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (mst_grp_6_wo_icb_rsp_ready               ),
  .o_icb_rsp_valid                (mst_grp_6_wo_icb_rsp_valid               ),
  .o_icb_rsp_err                  (mst_grp_6_wo_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (mst_grp_6_wo_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (mst_grp_6_wo_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (mst_grp_6_wo_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                slv_grp_0_icb_cmd_valid       ;
  wire                slv_grp_0_icb_cmd_ready       ;
  wire                slv_grp_0_icb_cmd_sel         ;
  wire                slv_grp_0_icb_cmd_read        ;
  wire    [  31:   0] slv_grp_0_icb_cmd_addr        ;
  wire    [  63:   0] slv_grp_0_icb_cmd_wdata       ;
  wire    [   7:   0] slv_grp_0_icb_cmd_wmask       ;
  wire    [   2:   0] slv_grp_0_icb_cmd_size        ;
  wire                slv_grp_0_icb_cmd_lock        ;
  wire                slv_grp_0_icb_cmd_excl        ;
  wire    [   7:   0] slv_grp_0_icb_cmd_xlen        ;
  wire    [   1:   0] slv_grp_0_icb_cmd_xburst      ;
  wire    [   1:   0] slv_grp_0_icb_cmd_modes       ;
  wire                slv_grp_0_icb_cmd_dmode       ;
  wire    [   2:   0] slv_grp_0_icb_cmd_attri       ;
  wire    [   1:   0] slv_grp_0_icb_cmd_beat        ;
  wire    [   2:   0] slv_grp_0_icb_cmd_usr         ;
  wire                slv_grp_0_icb_rsp_ready       ;
  wire                slv_grp_0_icb_rsp_valid       ;
  wire                slv_grp_0_icb_rsp_err         ;
  wire                slv_grp_0_icb_rsp_excl_ok     ;
  wire    [  63:   0] slv_grp_0_icb_rsp_rdata       ;
  wire    [   2:   0] slv_grp_0_icb_rsp_usr         ;
      wire                slv_grp_0_ro_icb_cmd_valid    ;
  wire                slv_grp_0_ro_icb_cmd_ready    ;
  wire                slv_grp_0_ro_icb_cmd_sel      ;
  wire                slv_grp_0_ro_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_0_ro_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_0_ro_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_0_ro_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_0_ro_icb_cmd_size     ;
  wire                slv_grp_0_ro_icb_cmd_lock     ;
  wire                slv_grp_0_ro_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_0_ro_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_0_ro_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_0_ro_icb_cmd_modes    ;
  wire                slv_grp_0_ro_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_0_ro_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_0_ro_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_0_ro_icb_cmd_usr      ;
  wire                slv_grp_0_ro_icb_rsp_ready    ;
  wire                slv_grp_0_ro_icb_rsp_valid    ;
  wire                slv_grp_0_ro_icb_rsp_err      ;
  wire                slv_grp_0_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_0_ro_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_0_ro_icb_rsp_usr      ;
      wire                slv_grp_0_wo_icb_cmd_valid    ;
  wire                slv_grp_0_wo_icb_cmd_ready    ;
  wire                slv_grp_0_wo_icb_cmd_sel      ;
  wire                slv_grp_0_wo_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_0_wo_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_0_wo_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_0_wo_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_0_wo_icb_cmd_size     ;
  wire                slv_grp_0_wo_icb_cmd_lock     ;
  wire                slv_grp_0_wo_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_0_wo_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_0_wo_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_0_wo_icb_cmd_modes    ;
  wire                slv_grp_0_wo_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_0_wo_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_0_wo_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_0_wo_icb_cmd_usr      ;
  wire                slv_grp_0_wo_icb_rsp_ready    ;
  wire                slv_grp_0_wo_icb_rsp_valid    ;
  wire                slv_grp_0_wo_icb_rsp_err      ;
  wire                slv_grp_0_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_0_wo_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_0_wo_icb_rsp_usr      ;
      wire                slv_grp0_p0_cmd_valid         ;
  wire                slv_grp0_p0_cmd_ready         ;
  wire                slv_grp0_p0_cmd_sel           ;
  wire                slv_grp0_p0_cmd_read          ;
  wire    [  31:   0] slv_grp0_p0_cmd_addr          ;
  wire    [  63:   0] slv_grp0_p0_cmd_wdata         ;
  wire    [   7:   0] slv_grp0_p0_cmd_wmask         ;
  wire    [   2:   0] slv_grp0_p0_cmd_size          ;
  wire                slv_grp0_p0_cmd_lock          ;
  wire                slv_grp0_p0_cmd_excl          ;
  wire    [   7:   0] slv_grp0_p0_cmd_xlen          ;
  wire    [   1:   0] slv_grp0_p0_cmd_xburst        ;
  wire    [   1:   0] slv_grp0_p0_cmd_modes         ;
  wire                slv_grp0_p0_cmd_dmode         ;
  wire    [   2:   0] slv_grp0_p0_cmd_attri         ;
  wire    [   1:   0] slv_grp0_p0_cmd_beat          ;
  wire    [   2:   0] slv_grp0_p0_cmd_usr           ;
  wire                slv_grp0_p0_rsp_ready         ;
  wire                slv_grp0_p0_rsp_valid         ;
  wire                slv_grp0_p0_rsp_err           ;
  wire                slv_grp0_p0_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp0_p0_rsp_rdata         ;
  wire    [   2:   0] slv_grp0_p0_rsp_usr           ;
      wire                slv_grp0_p0_w2n_cmd_valid     ;
  wire                slv_grp0_p0_w2n_cmd_ready     ;
  wire                slv_grp0_p0_w2n_cmd_sel       ;
  wire                slv_grp0_p0_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp0_p0_w2n_cmd_addr      ;
  wire    [  63:   0] slv_grp0_p0_w2n_cmd_wdata     ;
  wire    [   7:   0] slv_grp0_p0_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp0_p0_w2n_cmd_size      ;
  wire                slv_grp0_p0_w2n_cmd_lock      ;
  wire                slv_grp0_p0_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp0_p0_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp0_p0_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp0_p0_w2n_cmd_modes     ;
  wire                slv_grp0_p0_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp0_p0_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp0_p0_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp0_p0_w2n_cmd_usr       ;
  wire                slv_grp0_p0_w2n_rsp_ready     ;
  wire                slv_grp0_p0_w2n_rsp_valid     ;
  wire                slv_grp0_p0_w2n_rsp_err       ;
  wire                slv_grp0_p0_w2n_rsp_excl_ok   ;
  wire    [  63:   0] slv_grp0_p0_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp0_p0_w2n_rsp_usr       ;
      wire                slv_grp0_p0_ro_cmd_valid      ;
  wire                slv_grp0_p0_ro_cmd_ready      ;
  wire                slv_grp0_p0_ro_cmd_sel        ;
  wire                slv_grp0_p0_ro_cmd_read       ;
  wire    [  31:   0] slv_grp0_p0_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp0_p0_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp0_p0_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp0_p0_ro_cmd_size       ;
  wire                slv_grp0_p0_ro_cmd_lock       ;
  wire                slv_grp0_p0_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp0_p0_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp0_p0_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp0_p0_ro_cmd_modes      ;
  wire                slv_grp0_p0_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp0_p0_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp0_p0_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp0_p0_ro_cmd_usr        ;
  wire                slv_grp0_p0_ro_rsp_ready      ;
  wire                slv_grp0_p0_ro_rsp_valid      ;
  wire                slv_grp0_p0_ro_rsp_err        ;
  wire                slv_grp0_p0_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp0_p0_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp0_p0_ro_rsp_usr        ;
      wire                slv_grp0_p0_w2n_ro_cmd_valid  ;
  wire                slv_grp0_p0_w2n_ro_cmd_ready  ;
  wire                slv_grp0_p0_w2n_ro_cmd_sel    ;
  wire                slv_grp0_p0_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp0_p0_w2n_ro_cmd_addr   ;
  wire    [  63:   0] slv_grp0_p0_w2n_ro_cmd_wdata  ;
  wire    [   7:   0] slv_grp0_p0_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp0_p0_w2n_ro_cmd_size   ;
  wire                slv_grp0_p0_w2n_ro_cmd_lock   ;
  wire                slv_grp0_p0_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp0_p0_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp0_p0_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp0_p0_w2n_ro_cmd_modes  ;
  wire                slv_grp0_p0_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp0_p0_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp0_p0_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp0_p0_w2n_ro_cmd_usr    ;
  wire                slv_grp0_p0_w2n_ro_rsp_ready  ;
  wire                slv_grp0_p0_w2n_ro_rsp_valid  ;
  wire                slv_grp0_p0_w2n_ro_rsp_err    ;
  wire                slv_grp0_p0_w2n_ro_rsp_excl_ok ;
  wire    [  63:   0] slv_grp0_p0_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp0_p0_w2n_ro_rsp_usr    ;
      wire                slv_grp0_p0_wo_cmd_valid      ;
  wire                slv_grp0_p0_wo_cmd_ready      ;
  wire                slv_grp0_p0_wo_cmd_sel        ;
  wire                slv_grp0_p0_wo_cmd_read       ;
  wire    [  31:   0] slv_grp0_p0_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp0_p0_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp0_p0_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp0_p0_wo_cmd_size       ;
  wire                slv_grp0_p0_wo_cmd_lock       ;
  wire                slv_grp0_p0_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp0_p0_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp0_p0_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp0_p0_wo_cmd_modes      ;
  wire                slv_grp0_p0_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp0_p0_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp0_p0_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp0_p0_wo_cmd_usr        ;
  wire                slv_grp0_p0_wo_rsp_ready      ;
  wire                slv_grp0_p0_wo_rsp_valid      ;
  wire                slv_grp0_p0_wo_rsp_err        ;
  wire                slv_grp0_p0_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp0_p0_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp0_p0_wo_rsp_usr        ;
      wire                slv_grp0_p0_w2n_wo_cmd_valid  ;
  wire                slv_grp0_p0_w2n_wo_cmd_ready  ;
  wire                slv_grp0_p0_w2n_wo_cmd_sel    ;
  wire                slv_grp0_p0_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp0_p0_w2n_wo_cmd_addr   ;
  wire    [  63:   0] slv_grp0_p0_w2n_wo_cmd_wdata  ;
  wire    [   7:   0] slv_grp0_p0_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp0_p0_w2n_wo_cmd_size   ;
  wire                slv_grp0_p0_w2n_wo_cmd_lock   ;
  wire                slv_grp0_p0_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp0_p0_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp0_p0_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp0_p0_w2n_wo_cmd_modes  ;
  wire                slv_grp0_p0_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp0_p0_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp0_p0_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp0_p0_w2n_wo_cmd_usr    ;
  wire                slv_grp0_p0_w2n_wo_rsp_ready  ;
  wire                slv_grp0_p0_w2n_wo_rsp_valid  ;
  wire                slv_grp0_p0_w2n_wo_rsp_err    ;
  wire                slv_grp0_p0_w2n_wo_rsp_excl_ok ;
  wire    [  63:   0] slv_grp0_p0_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp0_p0_w2n_wo_rsp_usr    ;
                wire                      slv_grp0_p0_w2n_wo_rsp_last;
   e603_subsys_sgrp0_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1),
      .ICB_FIFO_CMD_DP        (1),
      .ICB_FIFO_RSP_DP        (0),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (32'h60000000),
      .O0_BASE_REGION_LSB(16),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (16 ),
      .SPLT_FIFO_OUTS_CNT_W(5),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp0_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_0_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (slv_grp_0_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (slv_grp_0_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (slv_grp_0_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (slv_grp_0_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_0_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_0_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_0_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_0_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (slv_grp_0_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (slv_grp_0_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_0_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_0_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_0_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (slv_grp_0_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_0_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_0_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_0_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (slv_grp_0_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (slv_grp_0_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (slv_grp_0_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (slv_grp_0_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_0_icb_rsp_usr         [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (slv_grp0_p0_cmd_valid                    ),
  .o0_icb_cmd_ready               (slv_grp0_p0_cmd_ready                    ),
  .o0_icb_cmd_sel                 (slv_grp0_p0_cmd_sel                      ),
  .o0_icb_cmd_read                (slv_grp0_p0_cmd_read                     ),
  .o0_icb_cmd_addr                (slv_grp0_p0_cmd_addr          [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp0_p0_cmd_wdata         [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp0_p0_cmd_wmask         [   7:   0]),
  .o0_icb_cmd_size                (slv_grp0_p0_cmd_size          [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp0_p0_cmd_lock                     ),
  .o0_icb_cmd_excl                (slv_grp0_p0_cmd_excl                     ),
  .o0_icb_cmd_xlen                (slv_grp0_p0_cmd_xlen          [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp0_p0_cmd_xburst        [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp0_p0_cmd_modes         [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp0_p0_cmd_dmode                    ),
  .o0_icb_cmd_attri               (slv_grp0_p0_cmd_attri         [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp0_p0_cmd_beat          [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp0_p0_cmd_usr           [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp0_p0_rsp_ready                    ),
  .o0_icb_rsp_valid               (slv_grp0_p0_rsp_valid                    ),
  .o0_icb_rsp_err                 (slv_grp0_p0_rsp_err                      ),
  .o0_icb_rsp_excl_ok             (slv_grp0_p0_rsp_excl_ok                  ),
  .o0_icb_rsp_rdata               (slv_grp0_p0_rsp_rdata         [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp0_p0_rsp_usr           [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (16),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_biu2iram_icb_icb_wconv(
        .i_icb_cmd_valid                (slv_grp0_p0_cmd_valid                    ),
  .i_icb_cmd_ready                (slv_grp0_p0_cmd_ready                    ),
  .i_icb_cmd_sel                  (slv_grp0_p0_cmd_sel                      ),
  .i_icb_cmd_read                 (slv_grp0_p0_cmd_read                     ),
  .i_icb_cmd_addr                 (slv_grp0_p0_cmd_addr          [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp0_p0_cmd_wdata         [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp0_p0_cmd_wmask         [   7:   0]),
  .i_icb_cmd_size                 (slv_grp0_p0_cmd_size          [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp0_p0_cmd_lock                     ),
  .i_icb_cmd_excl                 (slv_grp0_p0_cmd_excl                     ),
  .i_icb_cmd_xlen                 (slv_grp0_p0_cmd_xlen          [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp0_p0_cmd_xburst        [   1:   0]),
  .i_icb_cmd_modes                (slv_grp0_p0_cmd_modes         [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp0_p0_cmd_dmode                    ),
  .i_icb_cmd_attri                (slv_grp0_p0_cmd_attri         [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp0_p0_cmd_beat          [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp0_p0_cmd_usr           [   2:   0]),
  .i_icb_rsp_ready                (slv_grp0_p0_rsp_ready                    ),
  .i_icb_rsp_valid                (slv_grp0_p0_rsp_valid                    ),
  .i_icb_rsp_err                  (slv_grp0_p0_rsp_err                      ),
  .i_icb_rsp_excl_ok              (slv_grp0_p0_rsp_excl_ok                  ),
  .i_icb_rsp_rdata                (slv_grp0_p0_rsp_rdata         [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp0_p0_rsp_usr           [   2:   0]),
        .o_icb_cmd_valid                (slv_grp0_p0_w2n_cmd_valid                ),
  .o_icb_cmd_ready                (slv_grp0_p0_w2n_cmd_ready                ),
  .o_icb_cmd_sel                  (slv_grp0_p0_w2n_cmd_sel                  ),
  .o_icb_cmd_read                 (slv_grp0_p0_w2n_cmd_read                 ),
  .o_icb_cmd_addr                 (slv_grp0_p0_w2n_cmd_addr      [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp0_p0_w2n_cmd_wdata     [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp0_p0_w2n_cmd_wmask     [   7:   0]),
  .o_icb_cmd_size                 (slv_grp0_p0_w2n_cmd_size      [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp0_p0_w2n_cmd_lock                 ),
  .o_icb_cmd_excl                 (slv_grp0_p0_w2n_cmd_excl                 ),
  .o_icb_cmd_xlen                 (slv_grp0_p0_w2n_cmd_xlen      [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp0_p0_w2n_cmd_xburst    [   1:   0]),
  .o_icb_cmd_modes                (slv_grp0_p0_w2n_cmd_modes     [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp0_p0_w2n_cmd_dmode                ),
  .o_icb_cmd_attri                (slv_grp0_p0_w2n_cmd_attri     [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp0_p0_w2n_cmd_beat      [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp0_p0_w2n_cmd_usr       [   2:   0]),
  .o_icb_rsp_ready                (slv_grp0_p0_w2n_rsp_ready                ),
  .o_icb_rsp_valid                (slv_grp0_p0_w2n_rsp_valid                ),
  .o_icb_rsp_err                  (slv_grp0_p0_w2n_rsp_err                  ),
  .o_icb_rsp_excl_ok              (slv_grp0_p0_w2n_rsp_excl_ok              ),
  .o_icb_rsp_rdata                (slv_grp0_p0_w2n_rsp_rdata     [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp0_p0_w2n_rsp_usr       [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      assign slv_grp0_p0_w2n_rsp_usr = 3'b0;
      wire biu2iram_icb_bus_pend_active = 1'b0;
      wire biu2iram_icb_bus_icb_active;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(5+1)
      )u_biu2iram_icb__icb_active (
         .icb_active(biu2iram_icb_bus_icb_active),
            .icb_cmd_valid(slv_grp0_p0_w2n_cmd_valid),
            .icb_cmd_ready(slv_grp0_p0_w2n_cmd_ready),
            .icb_rsp_valid(slv_grp0_p0_w2n_rsp_valid),
            .icb_rsp_ready(slv_grp0_p0_w2n_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] biu2iram_icb_cmd_addr_full;
      assign biu2iram_icb_cmd_addr = biu2iram_icb_cmd_addr_full[16-1:0];
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(1),
    .O_SUPPORT_RATIO(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
    .OUTS_CNT_W   (5),
    .AW    (32),
    .DW    (64),
            .CMD_DP    (2),
            .RSP_DP    (2),
            .RSP_BYPBUF(0),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(0),
    .CMD_UW (1),
    .RSP_UW (1)
  )u_biu2iram_icb_icb_buffer(
    .i_clk_en (biu2iram_icb_clk_en),
    .o_clk_en (1'b1),
    .icb_buffer_active   (),
             .i_icb_cmd_usr(1'b0),
             .i_icb_rsp_usr(),
      .i_icb_cmd_valid                (slv_grp0_p0_w2n_cmd_valid                ),
  .i_icb_cmd_ready                (slv_grp0_p0_w2n_cmd_ready                ),
  .i_icb_cmd_sel                  (slv_grp0_p0_w2n_cmd_sel                  ),
  .i_icb_cmd_read                 (slv_grp0_p0_w2n_cmd_read                 ),
  .i_icb_cmd_addr                 (slv_grp0_p0_w2n_cmd_addr      [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp0_p0_w2n_cmd_wdata     [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp0_p0_w2n_cmd_wmask     [   7:   0]),
  .i_icb_cmd_size                 (slv_grp0_p0_w2n_cmd_size      [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp0_p0_w2n_cmd_lock                 ),
  .i_icb_cmd_excl                 (slv_grp0_p0_w2n_cmd_excl                 ),
  .i_icb_cmd_xlen                 (slv_grp0_p0_w2n_cmd_xlen      [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp0_p0_w2n_cmd_xburst    [   1:   0]),
  .i_icb_cmd_modes                (slv_grp0_p0_w2n_cmd_modes     [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp0_p0_w2n_cmd_dmode                ),
  .i_icb_cmd_attri                (slv_grp0_p0_w2n_cmd_attri     [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp0_p0_w2n_cmd_beat      [   1:   0]),
  .i_icb_rsp_ready                (slv_grp0_p0_w2n_rsp_ready                ),
  .i_icb_rsp_valid                (slv_grp0_p0_w2n_rsp_valid                ),
  .i_icb_rsp_err                  (slv_grp0_p0_w2n_rsp_err                  ),
  .i_icb_rsp_excl_ok              (slv_grp0_p0_w2n_rsp_excl_ok              ),
  .i_icb_rsp_rdata                (slv_grp0_p0_w2n_rsp_rdata     [  63:   0]),
      .o_icb_cmd_valid                (biu2iram_icb_cmd_valid                   ),
  .o_icb_cmd_ready                (biu2iram_icb_cmd_ready                   ),
  .o_icb_cmd_sel                  (biu2iram_icb_cmd_sel                     ),
  .o_icb_cmd_read                 (biu2iram_icb_cmd_read                    ),
  .o_icb_cmd_wdata                (biu2iram_icb_cmd_wdata        [  63:   0]),
  .o_icb_cmd_wmask                (biu2iram_icb_cmd_wmask        [   7:   0]),
  .o_icb_cmd_size                 (biu2iram_icb_cmd_size         [   2:   0]),
  .o_icb_cmd_lock                 (biu2iram_icb_cmd_lock                    ),
  .o_icb_cmd_excl                 (biu2iram_icb_cmd_excl                    ),
  .o_icb_cmd_xlen                 (biu2iram_icb_cmd_xlen         [   7:   0]),
  .o_icb_cmd_xburst               (biu2iram_icb_cmd_xburst       [   1:   0]),
  .o_icb_cmd_modes                (biu2iram_icb_cmd_modes        [   1:   0]),
  .o_icb_cmd_dmode                (biu2iram_icb_cmd_dmode                   ),
  .o_icb_cmd_attri                (biu2iram_icb_cmd_attri        [   2:   0]),
  .o_icb_cmd_beat                 (biu2iram_icb_cmd_beat         [   1:   0]),
  .o_icb_rsp_ready                (biu2iram_icb_rsp_ready                   ),
  .o_icb_rsp_valid                (biu2iram_icb_rsp_valid                   ),
  .o_icb_rsp_err                  (biu2iram_icb_rsp_err                     ),
  .o_icb_rsp_excl_ok              (biu2iram_icb_rsp_excl_ok                 ),
  .o_icb_rsp_rdata                (biu2iram_icb_rsp_rdata        [  63:   0]),
            .o_icb_cmd_usr(),
            .o_icb_rsp_usr(1'b0),
      .o_icb_cmd_addr(biu2iram_icb_cmd_addr_full),
      .clk  (biu2iram_icb_clk),
      .rst_n(biu2iram_icb_rst_n) 
  );
      wire                slv_grp_1_icb_cmd_valid       ;
  wire                slv_grp_1_icb_cmd_ready       ;
  wire                slv_grp_1_icb_cmd_sel         ;
  wire                slv_grp_1_icb_cmd_read        ;
  wire    [  31:   0] slv_grp_1_icb_cmd_addr        ;
  wire    [  63:   0] slv_grp_1_icb_cmd_wdata       ;
  wire    [   7:   0] slv_grp_1_icb_cmd_wmask       ;
  wire    [   2:   0] slv_grp_1_icb_cmd_size        ;
  wire                slv_grp_1_icb_cmd_lock        ;
  wire                slv_grp_1_icb_cmd_excl        ;
  wire    [   7:   0] slv_grp_1_icb_cmd_xlen        ;
  wire    [   1:   0] slv_grp_1_icb_cmd_xburst      ;
  wire    [   1:   0] slv_grp_1_icb_cmd_modes       ;
  wire                slv_grp_1_icb_cmd_dmode       ;
  wire    [   2:   0] slv_grp_1_icb_cmd_attri       ;
  wire    [   1:   0] slv_grp_1_icb_cmd_beat        ;
  wire    [   2:   0] slv_grp_1_icb_cmd_usr         ;
  wire                slv_grp_1_icb_rsp_ready       ;
  wire                slv_grp_1_icb_rsp_valid       ;
  wire                slv_grp_1_icb_rsp_err         ;
  wire                slv_grp_1_icb_rsp_excl_ok     ;
  wire    [  63:   0] slv_grp_1_icb_rsp_rdata       ;
  wire    [   2:   0] slv_grp_1_icb_rsp_usr         ;
      wire                slv_grp_1_ro_icb_cmd_valid    ;
  wire                slv_grp_1_ro_icb_cmd_ready    ;
  wire                slv_grp_1_ro_icb_cmd_sel      ;
  wire                slv_grp_1_ro_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_1_ro_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_1_ro_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_1_ro_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_1_ro_icb_cmd_size     ;
  wire                slv_grp_1_ro_icb_cmd_lock     ;
  wire                slv_grp_1_ro_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_1_ro_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_1_ro_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_1_ro_icb_cmd_modes    ;
  wire                slv_grp_1_ro_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_1_ro_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_1_ro_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_1_ro_icb_cmd_usr      ;
  wire                slv_grp_1_ro_icb_rsp_ready    ;
  wire                slv_grp_1_ro_icb_rsp_valid    ;
  wire                slv_grp_1_ro_icb_rsp_err      ;
  wire                slv_grp_1_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_1_ro_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_1_ro_icb_rsp_usr      ;
      wire                slv_grp_1_wo_icb_cmd_valid    ;
  wire                slv_grp_1_wo_icb_cmd_ready    ;
  wire                slv_grp_1_wo_icb_cmd_sel      ;
  wire                slv_grp_1_wo_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_1_wo_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_1_wo_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_1_wo_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_1_wo_icb_cmd_size     ;
  wire                slv_grp_1_wo_icb_cmd_lock     ;
  wire                slv_grp_1_wo_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_1_wo_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_1_wo_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_1_wo_icb_cmd_modes    ;
  wire                slv_grp_1_wo_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_1_wo_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_1_wo_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_1_wo_icb_cmd_usr      ;
  wire                slv_grp_1_wo_icb_rsp_ready    ;
  wire                slv_grp_1_wo_icb_rsp_valid    ;
  wire                slv_grp_1_wo_icb_rsp_err      ;
  wire                slv_grp_1_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_1_wo_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_1_wo_icb_rsp_usr      ;
      wire                slv_grp1_p0_cmd_valid         ;
  wire                slv_grp1_p0_cmd_ready         ;
  wire                slv_grp1_p0_cmd_sel           ;
  wire                slv_grp1_p0_cmd_read          ;
  wire    [  31:   0] slv_grp1_p0_cmd_addr          ;
  wire    [  63:   0] slv_grp1_p0_cmd_wdata         ;
  wire    [   7:   0] slv_grp1_p0_cmd_wmask         ;
  wire    [   2:   0] slv_grp1_p0_cmd_size          ;
  wire                slv_grp1_p0_cmd_lock          ;
  wire                slv_grp1_p0_cmd_excl          ;
  wire    [   7:   0] slv_grp1_p0_cmd_xlen          ;
  wire    [   1:   0] slv_grp1_p0_cmd_xburst        ;
  wire    [   1:   0] slv_grp1_p0_cmd_modes         ;
  wire                slv_grp1_p0_cmd_dmode         ;
  wire    [   2:   0] slv_grp1_p0_cmd_attri         ;
  wire    [   1:   0] slv_grp1_p0_cmd_beat          ;
  wire    [   2:   0] slv_grp1_p0_cmd_usr           ;
  wire                slv_grp1_p0_rsp_ready         ;
  wire                slv_grp1_p0_rsp_valid         ;
  wire                slv_grp1_p0_rsp_err           ;
  wire                slv_grp1_p0_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp1_p0_rsp_rdata         ;
  wire    [   2:   0] slv_grp1_p0_rsp_usr           ;
      wire                slv_grp1_p0_w2n_cmd_valid     ;
  wire                slv_grp1_p0_w2n_cmd_ready     ;
  wire                slv_grp1_p0_w2n_cmd_sel       ;
  wire                slv_grp1_p0_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp1_p0_w2n_cmd_addr      ;
  wire    [  63:   0] slv_grp1_p0_w2n_cmd_wdata     ;
  wire    [   7:   0] slv_grp1_p0_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp1_p0_w2n_cmd_size      ;
  wire                slv_grp1_p0_w2n_cmd_lock      ;
  wire                slv_grp1_p0_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp1_p0_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp1_p0_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp1_p0_w2n_cmd_modes     ;
  wire                slv_grp1_p0_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp1_p0_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp1_p0_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp1_p0_w2n_cmd_usr       ;
  wire                slv_grp1_p0_w2n_rsp_ready     ;
  wire                slv_grp1_p0_w2n_rsp_valid     ;
  wire                slv_grp1_p0_w2n_rsp_err       ;
  wire                slv_grp1_p0_w2n_rsp_excl_ok   ;
  wire    [  63:   0] slv_grp1_p0_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp1_p0_w2n_rsp_usr       ;
      wire                slv_grp1_p0_ro_cmd_valid      ;
  wire                slv_grp1_p0_ro_cmd_ready      ;
  wire                slv_grp1_p0_ro_cmd_sel        ;
  wire                slv_grp1_p0_ro_cmd_read       ;
  wire    [  31:   0] slv_grp1_p0_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp1_p0_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp1_p0_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp1_p0_ro_cmd_size       ;
  wire                slv_grp1_p0_ro_cmd_lock       ;
  wire                slv_grp1_p0_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp1_p0_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp1_p0_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp1_p0_ro_cmd_modes      ;
  wire                slv_grp1_p0_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp1_p0_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp1_p0_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp1_p0_ro_cmd_usr        ;
  wire                slv_grp1_p0_ro_rsp_ready      ;
  wire                slv_grp1_p0_ro_rsp_valid      ;
  wire                slv_grp1_p0_ro_rsp_err        ;
  wire                slv_grp1_p0_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp1_p0_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp1_p0_ro_rsp_usr        ;
      wire                slv_grp1_p0_w2n_ro_cmd_valid  ;
  wire                slv_grp1_p0_w2n_ro_cmd_ready  ;
  wire                slv_grp1_p0_w2n_ro_cmd_sel    ;
  wire                slv_grp1_p0_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp1_p0_w2n_ro_cmd_addr   ;
  wire    [  63:   0] slv_grp1_p0_w2n_ro_cmd_wdata  ;
  wire    [   7:   0] slv_grp1_p0_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp1_p0_w2n_ro_cmd_size   ;
  wire                slv_grp1_p0_w2n_ro_cmd_lock   ;
  wire                slv_grp1_p0_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp1_p0_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp1_p0_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp1_p0_w2n_ro_cmd_modes  ;
  wire                slv_grp1_p0_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp1_p0_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp1_p0_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp1_p0_w2n_ro_cmd_usr    ;
  wire                slv_grp1_p0_w2n_ro_rsp_ready  ;
  wire                slv_grp1_p0_w2n_ro_rsp_valid  ;
  wire                slv_grp1_p0_w2n_ro_rsp_err    ;
  wire                slv_grp1_p0_w2n_ro_rsp_excl_ok ;
  wire    [  63:   0] slv_grp1_p0_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp1_p0_w2n_ro_rsp_usr    ;
      wire                slv_grp1_p0_wo_cmd_valid      ;
  wire                slv_grp1_p0_wo_cmd_ready      ;
  wire                slv_grp1_p0_wo_cmd_sel        ;
  wire                slv_grp1_p0_wo_cmd_read       ;
  wire    [  31:   0] slv_grp1_p0_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp1_p0_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp1_p0_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp1_p0_wo_cmd_size       ;
  wire                slv_grp1_p0_wo_cmd_lock       ;
  wire                slv_grp1_p0_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp1_p0_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp1_p0_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp1_p0_wo_cmd_modes      ;
  wire                slv_grp1_p0_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp1_p0_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp1_p0_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp1_p0_wo_cmd_usr        ;
  wire                slv_grp1_p0_wo_rsp_ready      ;
  wire                slv_grp1_p0_wo_rsp_valid      ;
  wire                slv_grp1_p0_wo_rsp_err        ;
  wire                slv_grp1_p0_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp1_p0_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp1_p0_wo_rsp_usr        ;
      wire                slv_grp1_p0_w2n_wo_cmd_valid  ;
  wire                slv_grp1_p0_w2n_wo_cmd_ready  ;
  wire                slv_grp1_p0_w2n_wo_cmd_sel    ;
  wire                slv_grp1_p0_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp1_p0_w2n_wo_cmd_addr   ;
  wire    [  63:   0] slv_grp1_p0_w2n_wo_cmd_wdata  ;
  wire    [   7:   0] slv_grp1_p0_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp1_p0_w2n_wo_cmd_size   ;
  wire                slv_grp1_p0_w2n_wo_cmd_lock   ;
  wire                slv_grp1_p0_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp1_p0_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp1_p0_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp1_p0_w2n_wo_cmd_modes  ;
  wire                slv_grp1_p0_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp1_p0_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp1_p0_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp1_p0_w2n_wo_cmd_usr    ;
  wire                slv_grp1_p0_w2n_wo_rsp_ready  ;
  wire                slv_grp1_p0_w2n_wo_rsp_valid  ;
  wire                slv_grp1_p0_w2n_wo_rsp_err    ;
  wire                slv_grp1_p0_w2n_wo_rsp_excl_ok ;
  wire    [  63:   0] slv_grp1_p0_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp1_p0_w2n_wo_rsp_usr    ;
                wire                      slv_grp1_p0_w2n_wo_rsp_last;
   e603_subsys_sgrp1_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1),
      .ICB_FIFO_CMD_DP        (1),
      .ICB_FIFO_RSP_DP        (0),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (32'h68000000),
      .O0_BASE_REGION_LSB(16),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (16 ),
      .SPLT_FIFO_OUTS_CNT_W(5),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp1_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_1_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (slv_grp_1_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (slv_grp_1_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (slv_grp_1_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (slv_grp_1_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_1_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_1_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_1_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_1_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (slv_grp_1_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (slv_grp_1_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_1_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_1_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_1_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (slv_grp_1_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_1_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_1_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_1_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (slv_grp_1_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (slv_grp_1_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (slv_grp_1_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (slv_grp_1_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_1_icb_rsp_usr         [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (slv_grp1_p0_cmd_valid                    ),
  .o0_icb_cmd_ready               (slv_grp1_p0_cmd_ready                    ),
  .o0_icb_cmd_sel                 (slv_grp1_p0_cmd_sel                      ),
  .o0_icb_cmd_read                (slv_grp1_p0_cmd_read                     ),
  .o0_icb_cmd_addr                (slv_grp1_p0_cmd_addr          [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp1_p0_cmd_wdata         [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp1_p0_cmd_wmask         [   7:   0]),
  .o0_icb_cmd_size                (slv_grp1_p0_cmd_size          [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp1_p0_cmd_lock                     ),
  .o0_icb_cmd_excl                (slv_grp1_p0_cmd_excl                     ),
  .o0_icb_cmd_xlen                (slv_grp1_p0_cmd_xlen          [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp1_p0_cmd_xburst        [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp1_p0_cmd_modes         [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp1_p0_cmd_dmode                    ),
  .o0_icb_cmd_attri               (slv_grp1_p0_cmd_attri         [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp1_p0_cmd_beat          [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp1_p0_cmd_usr           [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp1_p0_rsp_ready                    ),
  .o0_icb_rsp_valid               (slv_grp1_p0_rsp_valid                    ),
  .o0_icb_rsp_err                 (slv_grp1_p0_rsp_err                      ),
  .o0_icb_rsp_excl_ok             (slv_grp1_p0_rsp_excl_ok                  ),
  .o0_icb_rsp_rdata               (slv_grp1_p0_rsp_rdata         [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp1_p0_rsp_usr           [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (16),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_biu2dram_icb_icb_wconv(
        .i_icb_cmd_valid                (slv_grp1_p0_cmd_valid                    ),
  .i_icb_cmd_ready                (slv_grp1_p0_cmd_ready                    ),
  .i_icb_cmd_sel                  (slv_grp1_p0_cmd_sel                      ),
  .i_icb_cmd_read                 (slv_grp1_p0_cmd_read                     ),
  .i_icb_cmd_addr                 (slv_grp1_p0_cmd_addr          [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp1_p0_cmd_wdata         [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp1_p0_cmd_wmask         [   7:   0]),
  .i_icb_cmd_size                 (slv_grp1_p0_cmd_size          [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp1_p0_cmd_lock                     ),
  .i_icb_cmd_excl                 (slv_grp1_p0_cmd_excl                     ),
  .i_icb_cmd_xlen                 (slv_grp1_p0_cmd_xlen          [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp1_p0_cmd_xburst        [   1:   0]),
  .i_icb_cmd_modes                (slv_grp1_p0_cmd_modes         [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp1_p0_cmd_dmode                    ),
  .i_icb_cmd_attri                (slv_grp1_p0_cmd_attri         [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp1_p0_cmd_beat          [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp1_p0_cmd_usr           [   2:   0]),
  .i_icb_rsp_ready                (slv_grp1_p0_rsp_ready                    ),
  .i_icb_rsp_valid                (slv_grp1_p0_rsp_valid                    ),
  .i_icb_rsp_err                  (slv_grp1_p0_rsp_err                      ),
  .i_icb_rsp_excl_ok              (slv_grp1_p0_rsp_excl_ok                  ),
  .i_icb_rsp_rdata                (slv_grp1_p0_rsp_rdata         [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp1_p0_rsp_usr           [   2:   0]),
        .o_icb_cmd_valid                (slv_grp1_p0_w2n_cmd_valid                ),
  .o_icb_cmd_ready                (slv_grp1_p0_w2n_cmd_ready                ),
  .o_icb_cmd_sel                  (slv_grp1_p0_w2n_cmd_sel                  ),
  .o_icb_cmd_read                 (slv_grp1_p0_w2n_cmd_read                 ),
  .o_icb_cmd_addr                 (slv_grp1_p0_w2n_cmd_addr      [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp1_p0_w2n_cmd_wdata     [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp1_p0_w2n_cmd_wmask     [   7:   0]),
  .o_icb_cmd_size                 (slv_grp1_p0_w2n_cmd_size      [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp1_p0_w2n_cmd_lock                 ),
  .o_icb_cmd_excl                 (slv_grp1_p0_w2n_cmd_excl                 ),
  .o_icb_cmd_xlen                 (slv_grp1_p0_w2n_cmd_xlen      [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp1_p0_w2n_cmd_xburst    [   1:   0]),
  .o_icb_cmd_modes                (slv_grp1_p0_w2n_cmd_modes     [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp1_p0_w2n_cmd_dmode                ),
  .o_icb_cmd_attri                (slv_grp1_p0_w2n_cmd_attri     [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp1_p0_w2n_cmd_beat      [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp1_p0_w2n_cmd_usr       [   2:   0]),
  .o_icb_rsp_ready                (slv_grp1_p0_w2n_rsp_ready                ),
  .o_icb_rsp_valid                (slv_grp1_p0_w2n_rsp_valid                ),
  .o_icb_rsp_err                  (slv_grp1_p0_w2n_rsp_err                  ),
  .o_icb_rsp_excl_ok              (slv_grp1_p0_w2n_rsp_excl_ok              ),
  .o_icb_rsp_rdata                (slv_grp1_p0_w2n_rsp_rdata     [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp1_p0_w2n_rsp_usr       [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      assign slv_grp1_p0_w2n_rsp_usr = 3'b0;
      wire biu2dram_icb_bus_pend_active = 1'b0;
      wire biu2dram_icb_bus_icb_active;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(5+1)
      )u_biu2dram_icb__icb_active (
         .icb_active(biu2dram_icb_bus_icb_active),
            .icb_cmd_valid(slv_grp1_p0_w2n_cmd_valid),
            .icb_cmd_ready(slv_grp1_p0_w2n_cmd_ready),
            .icb_rsp_valid(slv_grp1_p0_w2n_rsp_valid),
            .icb_rsp_ready(slv_grp1_p0_w2n_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] biu2dram_icb_cmd_addr_full;
      assign biu2dram_icb_cmd_addr = biu2dram_icb_cmd_addr_full[16-1:0];
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(1),
    .O_SUPPORT_RATIO(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
    .OUTS_CNT_W   (5),
    .AW    (32),
    .DW    (64),
            .CMD_DP    (2),
            .RSP_DP    (2),
            .RSP_BYPBUF(0),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(0),
    .CMD_UW (1),
    .RSP_UW (1)
  )u_biu2dram_icb_icb_buffer(
    .i_clk_en (biu2dram_icb_clk_en),
    .o_clk_en (1'b1),
    .icb_buffer_active   (),
             .i_icb_cmd_usr(1'b0),
             .i_icb_rsp_usr(),
      .i_icb_cmd_valid                (slv_grp1_p0_w2n_cmd_valid                ),
  .i_icb_cmd_ready                (slv_grp1_p0_w2n_cmd_ready                ),
  .i_icb_cmd_sel                  (slv_grp1_p0_w2n_cmd_sel                  ),
  .i_icb_cmd_read                 (slv_grp1_p0_w2n_cmd_read                 ),
  .i_icb_cmd_addr                 (slv_grp1_p0_w2n_cmd_addr      [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp1_p0_w2n_cmd_wdata     [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp1_p0_w2n_cmd_wmask     [   7:   0]),
  .i_icb_cmd_size                 (slv_grp1_p0_w2n_cmd_size      [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp1_p0_w2n_cmd_lock                 ),
  .i_icb_cmd_excl                 (slv_grp1_p0_w2n_cmd_excl                 ),
  .i_icb_cmd_xlen                 (slv_grp1_p0_w2n_cmd_xlen      [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp1_p0_w2n_cmd_xburst    [   1:   0]),
  .i_icb_cmd_modes                (slv_grp1_p0_w2n_cmd_modes     [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp1_p0_w2n_cmd_dmode                ),
  .i_icb_cmd_attri                (slv_grp1_p0_w2n_cmd_attri     [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp1_p0_w2n_cmd_beat      [   1:   0]),
  .i_icb_rsp_ready                (slv_grp1_p0_w2n_rsp_ready                ),
  .i_icb_rsp_valid                (slv_grp1_p0_w2n_rsp_valid                ),
  .i_icb_rsp_err                  (slv_grp1_p0_w2n_rsp_err                  ),
  .i_icb_rsp_excl_ok              (slv_grp1_p0_w2n_rsp_excl_ok              ),
  .i_icb_rsp_rdata                (slv_grp1_p0_w2n_rsp_rdata     [  63:   0]),
      .o_icb_cmd_valid                (biu2dram_icb_cmd_valid                   ),
  .o_icb_cmd_ready                (biu2dram_icb_cmd_ready                   ),
  .o_icb_cmd_sel                  (biu2dram_icb_cmd_sel                     ),
  .o_icb_cmd_read                 (biu2dram_icb_cmd_read                    ),
  .o_icb_cmd_wdata                (biu2dram_icb_cmd_wdata        [  63:   0]),
  .o_icb_cmd_wmask                (biu2dram_icb_cmd_wmask        [   7:   0]),
  .o_icb_cmd_size                 (biu2dram_icb_cmd_size         [   2:   0]),
  .o_icb_cmd_lock                 (biu2dram_icb_cmd_lock                    ),
  .o_icb_cmd_excl                 (biu2dram_icb_cmd_excl                    ),
  .o_icb_cmd_xlen                 (biu2dram_icb_cmd_xlen         [   7:   0]),
  .o_icb_cmd_xburst               (biu2dram_icb_cmd_xburst       [   1:   0]),
  .o_icb_cmd_modes                (biu2dram_icb_cmd_modes        [   1:   0]),
  .o_icb_cmd_dmode                (biu2dram_icb_cmd_dmode                   ),
  .o_icb_cmd_attri                (biu2dram_icb_cmd_attri        [   2:   0]),
  .o_icb_cmd_beat                 (biu2dram_icb_cmd_beat         [   1:   0]),
  .o_icb_rsp_ready                (biu2dram_icb_rsp_ready                   ),
  .o_icb_rsp_valid                (biu2dram_icb_rsp_valid                   ),
  .o_icb_rsp_err                  (biu2dram_icb_rsp_err                     ),
  .o_icb_rsp_excl_ok              (biu2dram_icb_rsp_excl_ok                 ),
  .o_icb_rsp_rdata                (biu2dram_icb_rsp_rdata        [  63:   0]),
            .o_icb_cmd_usr(),
            .o_icb_rsp_usr(1'b0),
      .o_icb_cmd_addr(biu2dram_icb_cmd_addr_full),
      .clk  (biu2dram_icb_clk),
      .rst_n(biu2dram_icb_rst_n) 
  );
      wire                slv_grp_2_icb_cmd_valid       ;
  wire                slv_grp_2_icb_cmd_ready       ;
  wire                slv_grp_2_icb_cmd_sel         ;
  wire                slv_grp_2_icb_cmd_read        ;
  wire    [  31:   0] slv_grp_2_icb_cmd_addr        ;
  wire    [  63:   0] slv_grp_2_icb_cmd_wdata       ;
  wire    [   7:   0] slv_grp_2_icb_cmd_wmask       ;
  wire    [   2:   0] slv_grp_2_icb_cmd_size        ;
  wire                slv_grp_2_icb_cmd_lock        ;
  wire                slv_grp_2_icb_cmd_excl        ;
  wire    [   7:   0] slv_grp_2_icb_cmd_xlen        ;
  wire    [   1:   0] slv_grp_2_icb_cmd_xburst      ;
  wire    [   1:   0] slv_grp_2_icb_cmd_modes       ;
  wire                slv_grp_2_icb_cmd_dmode       ;
  wire    [   2:   0] slv_grp_2_icb_cmd_attri       ;
  wire    [   1:   0] slv_grp_2_icb_cmd_beat        ;
  wire    [   2:   0] slv_grp_2_icb_cmd_usr         ;
  wire                slv_grp_2_icb_rsp_ready       ;
  wire                slv_grp_2_icb_rsp_valid       ;
  wire                slv_grp_2_icb_rsp_err         ;
  wire                slv_grp_2_icb_rsp_excl_ok     ;
  wire    [  63:   0] slv_grp_2_icb_rsp_rdata       ;
  wire    [   2:   0] slv_grp_2_icb_rsp_usr         ;
      wire                slv_grp_2_ro_icb_cmd_valid    ;
  wire                slv_grp_2_ro_icb_cmd_ready    ;
  wire                slv_grp_2_ro_icb_cmd_sel      ;
  wire                slv_grp_2_ro_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_2_ro_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_2_ro_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_2_ro_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_2_ro_icb_cmd_size     ;
  wire                slv_grp_2_ro_icb_cmd_lock     ;
  wire                slv_grp_2_ro_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_2_ro_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_2_ro_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_2_ro_icb_cmd_modes    ;
  wire                slv_grp_2_ro_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_2_ro_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_2_ro_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_2_ro_icb_cmd_usr      ;
  wire                slv_grp_2_ro_icb_rsp_ready    ;
  wire                slv_grp_2_ro_icb_rsp_valid    ;
  wire                slv_grp_2_ro_icb_rsp_err      ;
  wire                slv_grp_2_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_2_ro_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_2_ro_icb_rsp_usr      ;
      wire                slv_grp_2_wo_icb_cmd_valid    ;
  wire                slv_grp_2_wo_icb_cmd_ready    ;
  wire                slv_grp_2_wo_icb_cmd_sel      ;
  wire                slv_grp_2_wo_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_2_wo_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_2_wo_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_2_wo_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_2_wo_icb_cmd_size     ;
  wire                slv_grp_2_wo_icb_cmd_lock     ;
  wire                slv_grp_2_wo_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_2_wo_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_2_wo_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_2_wo_icb_cmd_modes    ;
  wire                slv_grp_2_wo_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_2_wo_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_2_wo_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_2_wo_icb_cmd_usr      ;
  wire                slv_grp_2_wo_icb_rsp_ready    ;
  wire                slv_grp_2_wo_icb_rsp_valid    ;
  wire                slv_grp_2_wo_icb_rsp_err      ;
  wire                slv_grp_2_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_2_wo_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_2_wo_icb_rsp_usr      ;
      wire                slv_grp2_p0_cmd_valid         ;
  wire                slv_grp2_p0_cmd_ready         ;
  wire                slv_grp2_p0_cmd_sel           ;
  wire                slv_grp2_p0_cmd_read          ;
  wire    [  31:   0] slv_grp2_p0_cmd_addr          ;
  wire    [  63:   0] slv_grp2_p0_cmd_wdata         ;
  wire    [   7:   0] slv_grp2_p0_cmd_wmask         ;
  wire    [   2:   0] slv_grp2_p0_cmd_size          ;
  wire                slv_grp2_p0_cmd_lock          ;
  wire                slv_grp2_p0_cmd_excl          ;
  wire    [   7:   0] slv_grp2_p0_cmd_xlen          ;
  wire    [   1:   0] slv_grp2_p0_cmd_xburst        ;
  wire    [   1:   0] slv_grp2_p0_cmd_modes         ;
  wire                slv_grp2_p0_cmd_dmode         ;
  wire    [   2:   0] slv_grp2_p0_cmd_attri         ;
  wire    [   1:   0] slv_grp2_p0_cmd_beat          ;
  wire    [   2:   0] slv_grp2_p0_cmd_usr           ;
  wire                slv_grp2_p0_rsp_ready         ;
  wire                slv_grp2_p0_rsp_valid         ;
  wire                slv_grp2_p0_rsp_err           ;
  wire                slv_grp2_p0_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp2_p0_rsp_rdata         ;
  wire    [   2:   0] slv_grp2_p0_rsp_usr           ;
      wire                slv_grp2_p0_w2n_cmd_valid     ;
  wire                slv_grp2_p0_w2n_cmd_ready     ;
  wire                slv_grp2_p0_w2n_cmd_sel       ;
  wire                slv_grp2_p0_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp2_p0_w2n_cmd_addr      ;
  wire    [  31:   0] slv_grp2_p0_w2n_cmd_wdata     ;
  wire    [   3:   0] slv_grp2_p0_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp2_p0_w2n_cmd_size      ;
  wire                slv_grp2_p0_w2n_cmd_lock      ;
  wire                slv_grp2_p0_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp2_p0_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp2_p0_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp2_p0_w2n_cmd_modes     ;
  wire                slv_grp2_p0_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp2_p0_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp2_p0_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp2_p0_w2n_cmd_usr       ;
  wire                slv_grp2_p0_w2n_rsp_ready     ;
  wire                slv_grp2_p0_w2n_rsp_valid     ;
  wire                slv_grp2_p0_w2n_rsp_err       ;
  wire                slv_grp2_p0_w2n_rsp_excl_ok   ;
  wire    [  31:   0] slv_grp2_p0_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp2_p0_w2n_rsp_usr       ;
      wire                slv_grp2_p0_ro_cmd_valid      ;
  wire                slv_grp2_p0_ro_cmd_ready      ;
  wire                slv_grp2_p0_ro_cmd_sel        ;
  wire                slv_grp2_p0_ro_cmd_read       ;
  wire    [  31:   0] slv_grp2_p0_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp2_p0_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp2_p0_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp2_p0_ro_cmd_size       ;
  wire                slv_grp2_p0_ro_cmd_lock       ;
  wire                slv_grp2_p0_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp2_p0_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp2_p0_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp2_p0_ro_cmd_modes      ;
  wire                slv_grp2_p0_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp2_p0_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp2_p0_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp2_p0_ro_cmd_usr        ;
  wire                slv_grp2_p0_ro_rsp_ready      ;
  wire                slv_grp2_p0_ro_rsp_valid      ;
  wire                slv_grp2_p0_ro_rsp_err        ;
  wire                slv_grp2_p0_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp2_p0_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp2_p0_ro_rsp_usr        ;
      wire                slv_grp2_p0_w2n_ro_cmd_valid  ;
  wire                slv_grp2_p0_w2n_ro_cmd_ready  ;
  wire                slv_grp2_p0_w2n_ro_cmd_sel    ;
  wire                slv_grp2_p0_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp2_p0_w2n_ro_cmd_addr   ;
  wire    [  31:   0] slv_grp2_p0_w2n_ro_cmd_wdata  ;
  wire    [   3:   0] slv_grp2_p0_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp2_p0_w2n_ro_cmd_size   ;
  wire                slv_grp2_p0_w2n_ro_cmd_lock   ;
  wire                slv_grp2_p0_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp2_p0_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp2_p0_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp2_p0_w2n_ro_cmd_modes  ;
  wire                slv_grp2_p0_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp2_p0_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp2_p0_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp2_p0_w2n_ro_cmd_usr    ;
  wire                slv_grp2_p0_w2n_ro_rsp_ready  ;
  wire                slv_grp2_p0_w2n_ro_rsp_valid  ;
  wire                slv_grp2_p0_w2n_ro_rsp_err    ;
  wire                slv_grp2_p0_w2n_ro_rsp_excl_ok ;
  wire    [  31:   0] slv_grp2_p0_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp2_p0_w2n_ro_rsp_usr    ;
      wire                slv_grp2_p0_wo_cmd_valid      ;
  wire                slv_grp2_p0_wo_cmd_ready      ;
  wire                slv_grp2_p0_wo_cmd_sel        ;
  wire                slv_grp2_p0_wo_cmd_read       ;
  wire    [  31:   0] slv_grp2_p0_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp2_p0_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp2_p0_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp2_p0_wo_cmd_size       ;
  wire                slv_grp2_p0_wo_cmd_lock       ;
  wire                slv_grp2_p0_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp2_p0_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp2_p0_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp2_p0_wo_cmd_modes      ;
  wire                slv_grp2_p0_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp2_p0_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp2_p0_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp2_p0_wo_cmd_usr        ;
  wire                slv_grp2_p0_wo_rsp_ready      ;
  wire                slv_grp2_p0_wo_rsp_valid      ;
  wire                slv_grp2_p0_wo_rsp_err        ;
  wire                slv_grp2_p0_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp2_p0_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp2_p0_wo_rsp_usr        ;
      wire                slv_grp2_p0_w2n_wo_cmd_valid  ;
  wire                slv_grp2_p0_w2n_wo_cmd_ready  ;
  wire                slv_grp2_p0_w2n_wo_cmd_sel    ;
  wire                slv_grp2_p0_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp2_p0_w2n_wo_cmd_addr   ;
  wire    [  31:   0] slv_grp2_p0_w2n_wo_cmd_wdata  ;
  wire    [   3:   0] slv_grp2_p0_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp2_p0_w2n_wo_cmd_size   ;
  wire                slv_grp2_p0_w2n_wo_cmd_lock   ;
  wire                slv_grp2_p0_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp2_p0_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp2_p0_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp2_p0_w2n_wo_cmd_modes  ;
  wire                slv_grp2_p0_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp2_p0_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp2_p0_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp2_p0_w2n_wo_cmd_usr    ;
  wire                slv_grp2_p0_w2n_wo_rsp_ready  ;
  wire                slv_grp2_p0_w2n_wo_rsp_valid  ;
  wire                slv_grp2_p0_w2n_wo_rsp_err    ;
  wire                slv_grp2_p0_w2n_wo_rsp_excl_ok ;
  wire    [  31:   0] slv_grp2_p0_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp2_p0_w2n_wo_rsp_usr    ;
                wire                      slv_grp2_p0_w2n_wo_rsp_last;
   e603_subsys_sgrp2_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (0),
      .ICB_FIFO_CMD_DP        (8),
      .ICB_FIFO_RSP_DP        (8),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (32'h0),
      .O0_BASE_REGION_LSB(12),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (16 ),
      .SPLT_FIFO_OUTS_CNT_W(5),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp2_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_2_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (slv_grp_2_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (slv_grp_2_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (slv_grp_2_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (slv_grp_2_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_2_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_2_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_2_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_2_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (slv_grp_2_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (slv_grp_2_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_2_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_2_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_2_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (slv_grp_2_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_2_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_2_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_2_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (slv_grp_2_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (slv_grp_2_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (slv_grp_2_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (slv_grp_2_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_2_icb_rsp_usr         [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (slv_grp2_p0_cmd_valid                    ),
  .o0_icb_cmd_ready               (slv_grp2_p0_cmd_ready                    ),
  .o0_icb_cmd_sel                 (slv_grp2_p0_cmd_sel                      ),
  .o0_icb_cmd_read                (slv_grp2_p0_cmd_read                     ),
  .o0_icb_cmd_addr                (slv_grp2_p0_cmd_addr          [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp2_p0_cmd_wdata         [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp2_p0_cmd_wmask         [   7:   0]),
  .o0_icb_cmd_size                (slv_grp2_p0_cmd_size          [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp2_p0_cmd_lock                     ),
  .o0_icb_cmd_excl                (slv_grp2_p0_cmd_excl                     ),
  .o0_icb_cmd_xlen                (slv_grp2_p0_cmd_xlen          [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp2_p0_cmd_xburst        [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp2_p0_cmd_modes         [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp2_p0_cmd_dmode                    ),
  .o0_icb_cmd_attri               (slv_grp2_p0_cmd_attri         [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp2_p0_cmd_beat          [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp2_p0_cmd_usr           [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp2_p0_rsp_ready                    ),
  .o0_icb_rsp_valid               (slv_grp2_p0_rsp_valid                    ),
  .o0_icb_rsp_err                 (slv_grp2_p0_rsp_err                      ),
  .o0_icb_rsp_excl_ok             (slv_grp2_p0_rsp_excl_ok                  ),
  .o0_icb_rsp_rdata               (slv_grp2_p0_rsp_rdata         [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp2_p0_rsp_usr           [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (16),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(32 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_addr0_icb_icb_wconv(
        .i_icb_cmd_valid                (slv_grp2_p0_cmd_valid                    ),
  .i_icb_cmd_ready                (slv_grp2_p0_cmd_ready                    ),
  .i_icb_cmd_sel                  (slv_grp2_p0_cmd_sel                      ),
  .i_icb_cmd_read                 (slv_grp2_p0_cmd_read                     ),
  .i_icb_cmd_addr                 (slv_grp2_p0_cmd_addr          [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp2_p0_cmd_wdata         [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp2_p0_cmd_wmask         [   7:   0]),
  .i_icb_cmd_size                 (slv_grp2_p0_cmd_size          [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp2_p0_cmd_lock                     ),
  .i_icb_cmd_excl                 (slv_grp2_p0_cmd_excl                     ),
  .i_icb_cmd_xlen                 (slv_grp2_p0_cmd_xlen          [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp2_p0_cmd_xburst        [   1:   0]),
  .i_icb_cmd_modes                (slv_grp2_p0_cmd_modes         [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp2_p0_cmd_dmode                    ),
  .i_icb_cmd_attri                (slv_grp2_p0_cmd_attri         [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp2_p0_cmd_beat          [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp2_p0_cmd_usr           [   2:   0]),
  .i_icb_rsp_ready                (slv_grp2_p0_rsp_ready                    ),
  .i_icb_rsp_valid                (slv_grp2_p0_rsp_valid                    ),
  .i_icb_rsp_err                  (slv_grp2_p0_rsp_err                      ),
  .i_icb_rsp_excl_ok              (slv_grp2_p0_rsp_excl_ok                  ),
  .i_icb_rsp_rdata                (slv_grp2_p0_rsp_rdata         [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp2_p0_rsp_usr           [   2:   0]),
        .o_icb_cmd_valid                (slv_grp2_p0_w2n_cmd_valid                ),
  .o_icb_cmd_ready                (slv_grp2_p0_w2n_cmd_ready                ),
  .o_icb_cmd_sel                  (slv_grp2_p0_w2n_cmd_sel                  ),
  .o_icb_cmd_read                 (slv_grp2_p0_w2n_cmd_read                 ),
  .o_icb_cmd_addr                 (slv_grp2_p0_w2n_cmd_addr      [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp2_p0_w2n_cmd_wdata     [  31:   0]),
  .o_icb_cmd_wmask                (slv_grp2_p0_w2n_cmd_wmask     [   3:   0]),
  .o_icb_cmd_size                 (slv_grp2_p0_w2n_cmd_size      [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp2_p0_w2n_cmd_lock                 ),
  .o_icb_cmd_excl                 (slv_grp2_p0_w2n_cmd_excl                 ),
  .o_icb_cmd_xlen                 (slv_grp2_p0_w2n_cmd_xlen      [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp2_p0_w2n_cmd_xburst    [   1:   0]),
  .o_icb_cmd_modes                (slv_grp2_p0_w2n_cmd_modes     [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp2_p0_w2n_cmd_dmode                ),
  .o_icb_cmd_attri                (slv_grp2_p0_w2n_cmd_attri     [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp2_p0_w2n_cmd_beat      [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp2_p0_w2n_cmd_usr       [   2:   0]),
  .o_icb_rsp_ready                (slv_grp2_p0_w2n_rsp_ready                ),
  .o_icb_rsp_valid                (slv_grp2_p0_w2n_rsp_valid                ),
  .o_icb_rsp_err                  (slv_grp2_p0_w2n_rsp_err                  ),
  .o_icb_rsp_excl_ok              (slv_grp2_p0_w2n_rsp_excl_ok              ),
  .o_icb_rsp_rdata                (slv_grp2_p0_w2n_rsp_rdata     [  31:   0]),
  .o_icb_rsp_usr                  (slv_grp2_p0_w2n_rsp_usr       [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      assign slv_grp2_p0_w2n_rsp_usr = 3'b0;
      wire addr0_icb_bus_pend_active = 1'b0;
      wire addr0_icb_bus_icb_active;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(5+1)
      )u_addr0_icb__icb_active (
         .icb_active(addr0_icb_bus_icb_active),
            .icb_cmd_valid(slv_grp2_p0_w2n_cmd_valid),
            .icb_cmd_ready(slv_grp2_p0_w2n_cmd_ready),
            .icb_rsp_valid(slv_grp2_p0_w2n_rsp_valid),
            .icb_rsp_ready(slv_grp2_p0_w2n_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] addr0_icb_cmd_addr_full;
      assign addr0_icb_cmd_addr = addr0_icb_cmd_addr_full[32-1:0];
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(0),
    .O_SUPPORT_RATIO(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
    .OUTS_CNT_W   (5),
    .AW    (32),
    .DW    (32),
            .CMD_DP    (1),
            .RSP_DP    (1),
            .RSP_BYPBUF(0),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(1),
    .CMD_UW (1),
    .RSP_UW (1)
  )u_addr0_icb_icb_buffer(
    .i_clk_en (1'b1),
    .o_clk_en (1'b1),
    .icb_buffer_active   (),
             .i_icb_cmd_usr(1'b0),
             .i_icb_rsp_usr(),
      .i_icb_cmd_valid                (slv_grp2_p0_w2n_cmd_valid                ),
  .i_icb_cmd_ready                (slv_grp2_p0_w2n_cmd_ready                ),
  .i_icb_cmd_sel                  (slv_grp2_p0_w2n_cmd_sel                  ),
  .i_icb_cmd_read                 (slv_grp2_p0_w2n_cmd_read                 ),
  .i_icb_cmd_addr                 (slv_grp2_p0_w2n_cmd_addr      [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp2_p0_w2n_cmd_wdata     [  31:   0]),
  .i_icb_cmd_wmask                (slv_grp2_p0_w2n_cmd_wmask     [   3:   0]),
  .i_icb_cmd_size                 (slv_grp2_p0_w2n_cmd_size      [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp2_p0_w2n_cmd_lock                 ),
  .i_icb_cmd_excl                 (slv_grp2_p0_w2n_cmd_excl                 ),
  .i_icb_cmd_xlen                 (slv_grp2_p0_w2n_cmd_xlen      [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp2_p0_w2n_cmd_xburst    [   1:   0]),
  .i_icb_cmd_modes                (slv_grp2_p0_w2n_cmd_modes     [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp2_p0_w2n_cmd_dmode                ),
  .i_icb_cmd_attri                (slv_grp2_p0_w2n_cmd_attri     [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp2_p0_w2n_cmd_beat      [   1:   0]),
  .i_icb_rsp_ready                (slv_grp2_p0_w2n_rsp_ready                ),
  .i_icb_rsp_valid                (slv_grp2_p0_w2n_rsp_valid                ),
  .i_icb_rsp_err                  (slv_grp2_p0_w2n_rsp_err                  ),
  .i_icb_rsp_excl_ok              (slv_grp2_p0_w2n_rsp_excl_ok              ),
  .i_icb_rsp_rdata                (slv_grp2_p0_w2n_rsp_rdata     [  31:   0]),
      .o_icb_cmd_valid                (addr0_icb_cmd_valid                      ),
  .o_icb_cmd_ready                (addr0_icb_cmd_ready                      ),
  .o_icb_cmd_sel                  (addr0_icb_cmd_sel                        ),
  .o_icb_cmd_read                 (addr0_icb_cmd_read                       ),
  .o_icb_cmd_wdata                (addr0_icb_cmd_wdata           [  31:   0]),
  .o_icb_cmd_wmask                (addr0_icb_cmd_wmask           [   3:   0]),
  .o_icb_cmd_size                 (addr0_icb_cmd_size            [   2:   0]),
  .o_icb_cmd_lock                 (addr0_icb_cmd_lock                       ),
  .o_icb_cmd_excl                 (addr0_icb_cmd_excl                       ),
  .o_icb_cmd_xlen                 (addr0_icb_cmd_xlen            [   7:   0]),
  .o_icb_cmd_xburst               (addr0_icb_cmd_xburst          [   1:   0]),
  .o_icb_cmd_modes                (addr0_icb_cmd_modes           [   1:   0]),
  .o_icb_cmd_dmode                (addr0_icb_cmd_dmode                      ),
  .o_icb_cmd_attri                (addr0_icb_cmd_attri           [   2:   0]),
  .o_icb_cmd_beat                 (addr0_icb_cmd_beat            [   1:   0]),
  .o_icb_rsp_ready                (addr0_icb_rsp_ready                      ),
  .o_icb_rsp_valid                (addr0_icb_rsp_valid                      ),
  .o_icb_rsp_err                  (addr0_icb_rsp_err                        ),
  .o_icb_rsp_excl_ok              (addr0_icb_rsp_excl_ok                    ),
  .o_icb_rsp_rdata                (addr0_icb_rsp_rdata           [  31:   0]),
            .o_icb_cmd_usr(),
            .o_icb_rsp_usr(1'b0),
      .o_icb_cmd_addr(addr0_icb_cmd_addr_full),
      .clk  (clk_fab),  
      .rst_n(rst_n)
  );
      wire                slv_grp_3_icb_cmd_valid       ;
  wire                slv_grp_3_icb_cmd_ready       ;
  wire                slv_grp_3_icb_cmd_sel         ;
  wire                slv_grp_3_icb_cmd_read        ;
  wire    [  31:   0] slv_grp_3_icb_cmd_addr        ;
  wire    [  63:   0] slv_grp_3_icb_cmd_wdata       ;
  wire    [   7:   0] slv_grp_3_icb_cmd_wmask       ;
  wire    [   2:   0] slv_grp_3_icb_cmd_size        ;
  wire                slv_grp_3_icb_cmd_lock        ;
  wire                slv_grp_3_icb_cmd_excl        ;
  wire    [   7:   0] slv_grp_3_icb_cmd_xlen        ;
  wire    [   1:   0] slv_grp_3_icb_cmd_xburst      ;
  wire    [   1:   0] slv_grp_3_icb_cmd_modes       ;
  wire                slv_grp_3_icb_cmd_dmode       ;
  wire    [   2:   0] slv_grp_3_icb_cmd_attri       ;
  wire    [   1:   0] slv_grp_3_icb_cmd_beat        ;
  wire    [   2:   0] slv_grp_3_icb_cmd_usr         ;
  wire                slv_grp_3_icb_rsp_ready       ;
  wire                slv_grp_3_icb_rsp_valid       ;
  wire                slv_grp_3_icb_rsp_err         ;
  wire                slv_grp_3_icb_rsp_excl_ok     ;
  wire    [  63:   0] slv_grp_3_icb_rsp_rdata       ;
  wire    [   2:   0] slv_grp_3_icb_rsp_usr         ;
      wire                slv_grp_3_ro_icb_cmd_valid    ;
  wire                slv_grp_3_ro_icb_cmd_ready    ;
  wire                slv_grp_3_ro_icb_cmd_sel      ;
  wire                slv_grp_3_ro_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_3_ro_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_3_ro_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_3_ro_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_3_ro_icb_cmd_size     ;
  wire                slv_grp_3_ro_icb_cmd_lock     ;
  wire                slv_grp_3_ro_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_3_ro_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_3_ro_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_3_ro_icb_cmd_modes    ;
  wire                slv_grp_3_ro_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_3_ro_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_3_ro_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_3_ro_icb_cmd_usr      ;
  wire                slv_grp_3_ro_icb_rsp_ready    ;
  wire                slv_grp_3_ro_icb_rsp_valid    ;
  wire                slv_grp_3_ro_icb_rsp_err      ;
  wire                slv_grp_3_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_3_ro_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_3_ro_icb_rsp_usr      ;
      wire                slv_grp_3_wo_icb_cmd_valid    ;
  wire                slv_grp_3_wo_icb_cmd_ready    ;
  wire                slv_grp_3_wo_icb_cmd_sel      ;
  wire                slv_grp_3_wo_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_3_wo_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_3_wo_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_3_wo_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_3_wo_icb_cmd_size     ;
  wire                slv_grp_3_wo_icb_cmd_lock     ;
  wire                slv_grp_3_wo_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_3_wo_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_3_wo_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_3_wo_icb_cmd_modes    ;
  wire                slv_grp_3_wo_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_3_wo_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_3_wo_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_3_wo_icb_cmd_usr      ;
  wire                slv_grp_3_wo_icb_rsp_ready    ;
  wire                slv_grp_3_wo_icb_rsp_valid    ;
  wire                slv_grp_3_wo_icb_rsp_err      ;
  wire                slv_grp_3_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_3_wo_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_3_wo_icb_rsp_usr      ;
      wire                slv_grp3_p0_cmd_valid         ;
  wire                slv_grp3_p0_cmd_ready         ;
  wire                slv_grp3_p0_cmd_sel           ;
  wire                slv_grp3_p0_cmd_read          ;
  wire    [  31:   0] slv_grp3_p0_cmd_addr          ;
  wire    [  63:   0] slv_grp3_p0_cmd_wdata         ;
  wire    [   7:   0] slv_grp3_p0_cmd_wmask         ;
  wire    [   2:   0] slv_grp3_p0_cmd_size          ;
  wire                slv_grp3_p0_cmd_lock          ;
  wire                slv_grp3_p0_cmd_excl          ;
  wire    [   7:   0] slv_grp3_p0_cmd_xlen          ;
  wire    [   1:   0] slv_grp3_p0_cmd_xburst        ;
  wire    [   1:   0] slv_grp3_p0_cmd_modes         ;
  wire                slv_grp3_p0_cmd_dmode         ;
  wire    [   2:   0] slv_grp3_p0_cmd_attri         ;
  wire    [   1:   0] slv_grp3_p0_cmd_beat          ;
  wire    [   2:   0] slv_grp3_p0_cmd_usr           ;
  wire                slv_grp3_p0_rsp_ready         ;
  wire                slv_grp3_p0_rsp_valid         ;
  wire                slv_grp3_p0_rsp_err           ;
  wire                slv_grp3_p0_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp3_p0_rsp_rdata         ;
  wire    [   2:   0] slv_grp3_p0_rsp_usr           ;
      wire                slv_grp3_p0_w2n_cmd_valid     ;
  wire                slv_grp3_p0_w2n_cmd_ready     ;
  wire                slv_grp3_p0_w2n_cmd_sel       ;
  wire                slv_grp3_p0_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp3_p0_w2n_cmd_addr      ;
  wire    [  31:   0] slv_grp3_p0_w2n_cmd_wdata     ;
  wire    [   3:   0] slv_grp3_p0_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp3_p0_w2n_cmd_size      ;
  wire                slv_grp3_p0_w2n_cmd_lock      ;
  wire                slv_grp3_p0_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp3_p0_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp3_p0_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp3_p0_w2n_cmd_modes     ;
  wire                slv_grp3_p0_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp3_p0_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp3_p0_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp3_p0_w2n_cmd_usr       ;
  wire                slv_grp3_p0_w2n_rsp_ready     ;
  wire                slv_grp3_p0_w2n_rsp_valid     ;
  wire                slv_grp3_p0_w2n_rsp_err       ;
  wire                slv_grp3_p0_w2n_rsp_excl_ok   ;
  wire    [  31:   0] slv_grp3_p0_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp3_p0_w2n_rsp_usr       ;
      wire                slv_grp3_p0_ro_cmd_valid      ;
  wire                slv_grp3_p0_ro_cmd_ready      ;
  wire                slv_grp3_p0_ro_cmd_sel        ;
  wire                slv_grp3_p0_ro_cmd_read       ;
  wire    [  31:   0] slv_grp3_p0_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp3_p0_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp3_p0_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp3_p0_ro_cmd_size       ;
  wire                slv_grp3_p0_ro_cmd_lock       ;
  wire                slv_grp3_p0_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp3_p0_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp3_p0_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp3_p0_ro_cmd_modes      ;
  wire                slv_grp3_p0_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp3_p0_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp3_p0_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp3_p0_ro_cmd_usr        ;
  wire                slv_grp3_p0_ro_rsp_ready      ;
  wire                slv_grp3_p0_ro_rsp_valid      ;
  wire                slv_grp3_p0_ro_rsp_err        ;
  wire                slv_grp3_p0_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp3_p0_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp3_p0_ro_rsp_usr        ;
      wire                slv_grp3_p0_w2n_ro_cmd_valid  ;
  wire                slv_grp3_p0_w2n_ro_cmd_ready  ;
  wire                slv_grp3_p0_w2n_ro_cmd_sel    ;
  wire                slv_grp3_p0_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp3_p0_w2n_ro_cmd_addr   ;
  wire    [  31:   0] slv_grp3_p0_w2n_ro_cmd_wdata  ;
  wire    [   3:   0] slv_grp3_p0_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp3_p0_w2n_ro_cmd_size   ;
  wire                slv_grp3_p0_w2n_ro_cmd_lock   ;
  wire                slv_grp3_p0_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp3_p0_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp3_p0_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp3_p0_w2n_ro_cmd_modes  ;
  wire                slv_grp3_p0_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp3_p0_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp3_p0_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp3_p0_w2n_ro_cmd_usr    ;
  wire                slv_grp3_p0_w2n_ro_rsp_ready  ;
  wire                slv_grp3_p0_w2n_ro_rsp_valid  ;
  wire                slv_grp3_p0_w2n_ro_rsp_err    ;
  wire                slv_grp3_p0_w2n_ro_rsp_excl_ok ;
  wire    [  31:   0] slv_grp3_p0_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp3_p0_w2n_ro_rsp_usr    ;
      wire                slv_grp3_p0_wo_cmd_valid      ;
  wire                slv_grp3_p0_wo_cmd_ready      ;
  wire                slv_grp3_p0_wo_cmd_sel        ;
  wire                slv_grp3_p0_wo_cmd_read       ;
  wire    [  31:   0] slv_grp3_p0_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp3_p0_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp3_p0_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp3_p0_wo_cmd_size       ;
  wire                slv_grp3_p0_wo_cmd_lock       ;
  wire                slv_grp3_p0_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp3_p0_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp3_p0_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp3_p0_wo_cmd_modes      ;
  wire                slv_grp3_p0_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp3_p0_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp3_p0_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp3_p0_wo_cmd_usr        ;
  wire                slv_grp3_p0_wo_rsp_ready      ;
  wire                slv_grp3_p0_wo_rsp_valid      ;
  wire                slv_grp3_p0_wo_rsp_err        ;
  wire                slv_grp3_p0_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp3_p0_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp3_p0_wo_rsp_usr        ;
      wire                slv_grp3_p0_w2n_wo_cmd_valid  ;
  wire                slv_grp3_p0_w2n_wo_cmd_ready  ;
  wire                slv_grp3_p0_w2n_wo_cmd_sel    ;
  wire                slv_grp3_p0_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp3_p0_w2n_wo_cmd_addr   ;
  wire    [  31:   0] slv_grp3_p0_w2n_wo_cmd_wdata  ;
  wire    [   3:   0] slv_grp3_p0_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp3_p0_w2n_wo_cmd_size   ;
  wire                slv_grp3_p0_w2n_wo_cmd_lock   ;
  wire                slv_grp3_p0_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp3_p0_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp3_p0_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp3_p0_w2n_wo_cmd_modes  ;
  wire                slv_grp3_p0_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp3_p0_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp3_p0_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp3_p0_w2n_wo_cmd_usr    ;
  wire                slv_grp3_p0_w2n_wo_rsp_ready  ;
  wire                slv_grp3_p0_w2n_wo_rsp_valid  ;
  wire                slv_grp3_p0_w2n_wo_rsp_err    ;
  wire                slv_grp3_p0_w2n_wo_rsp_excl_ok ;
  wire    [  31:   0] slv_grp3_p0_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp3_p0_w2n_wo_rsp_usr    ;
                wire                      slv_grp3_p0_w2n_wo_rsp_last;
   e603_subsys_sgrp3_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (0),
      .ICB_FIFO_CMD_DP        (8),
      .ICB_FIFO_RSP_DP        (8),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (32'h20000000),
      .O0_BASE_REGION_LSB(28),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (16 ),
      .SPLT_FIFO_OUTS_CNT_W(5),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp3_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_3_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (slv_grp_3_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (slv_grp_3_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (slv_grp_3_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (slv_grp_3_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_3_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_3_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_3_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_3_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (slv_grp_3_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (slv_grp_3_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_3_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_3_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_3_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (slv_grp_3_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_3_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_3_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_3_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (slv_grp_3_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (slv_grp_3_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (slv_grp_3_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (slv_grp_3_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_3_icb_rsp_usr         [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (slv_grp3_p0_cmd_valid                    ),
  .o0_icb_cmd_ready               (slv_grp3_p0_cmd_ready                    ),
  .o0_icb_cmd_sel                 (slv_grp3_p0_cmd_sel                      ),
  .o0_icb_cmd_read                (slv_grp3_p0_cmd_read                     ),
  .o0_icb_cmd_addr                (slv_grp3_p0_cmd_addr          [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp3_p0_cmd_wdata         [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp3_p0_cmd_wmask         [   7:   0]),
  .o0_icb_cmd_size                (slv_grp3_p0_cmd_size          [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp3_p0_cmd_lock                     ),
  .o0_icb_cmd_excl                (slv_grp3_p0_cmd_excl                     ),
  .o0_icb_cmd_xlen                (slv_grp3_p0_cmd_xlen          [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp3_p0_cmd_xburst        [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp3_p0_cmd_modes         [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp3_p0_cmd_dmode                    ),
  .o0_icb_cmd_attri               (slv_grp3_p0_cmd_attri         [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp3_p0_cmd_beat          [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp3_p0_cmd_usr           [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp3_p0_rsp_ready                    ),
  .o0_icb_rsp_valid               (slv_grp3_p0_rsp_valid                    ),
  .o0_icb_rsp_err                 (slv_grp3_p0_rsp_err                      ),
  .o0_icb_rsp_excl_ok             (slv_grp3_p0_rsp_excl_ok                  ),
  .o0_icb_rsp_rdata               (slv_grp3_p0_rsp_rdata         [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp3_p0_rsp_usr           [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (16),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(32 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_qspi0_ro_icb_icb_wconv(
        .i_icb_cmd_valid                (slv_grp3_p0_cmd_valid                    ),
  .i_icb_cmd_ready                (slv_grp3_p0_cmd_ready                    ),
  .i_icb_cmd_sel                  (slv_grp3_p0_cmd_sel                      ),
  .i_icb_cmd_read                 (slv_grp3_p0_cmd_read                     ),
  .i_icb_cmd_addr                 (slv_grp3_p0_cmd_addr          [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp3_p0_cmd_wdata         [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp3_p0_cmd_wmask         [   7:   0]),
  .i_icb_cmd_size                 (slv_grp3_p0_cmd_size          [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp3_p0_cmd_lock                     ),
  .i_icb_cmd_excl                 (slv_grp3_p0_cmd_excl                     ),
  .i_icb_cmd_xlen                 (slv_grp3_p0_cmd_xlen          [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp3_p0_cmd_xburst        [   1:   0]),
  .i_icb_cmd_modes                (slv_grp3_p0_cmd_modes         [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp3_p0_cmd_dmode                    ),
  .i_icb_cmd_attri                (slv_grp3_p0_cmd_attri         [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp3_p0_cmd_beat          [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp3_p0_cmd_usr           [   2:   0]),
  .i_icb_rsp_ready                (slv_grp3_p0_rsp_ready                    ),
  .i_icb_rsp_valid                (slv_grp3_p0_rsp_valid                    ),
  .i_icb_rsp_err                  (slv_grp3_p0_rsp_err                      ),
  .i_icb_rsp_excl_ok              (slv_grp3_p0_rsp_excl_ok                  ),
  .i_icb_rsp_rdata                (slv_grp3_p0_rsp_rdata         [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp3_p0_rsp_usr           [   2:   0]),
        .o_icb_cmd_valid                (slv_grp3_p0_w2n_cmd_valid                ),
  .o_icb_cmd_ready                (slv_grp3_p0_w2n_cmd_ready                ),
  .o_icb_cmd_sel                  (slv_grp3_p0_w2n_cmd_sel                  ),
  .o_icb_cmd_read                 (slv_grp3_p0_w2n_cmd_read                 ),
  .o_icb_cmd_addr                 (slv_grp3_p0_w2n_cmd_addr      [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp3_p0_w2n_cmd_wdata     [  31:   0]),
  .o_icb_cmd_wmask                (slv_grp3_p0_w2n_cmd_wmask     [   3:   0]),
  .o_icb_cmd_size                 (slv_grp3_p0_w2n_cmd_size      [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp3_p0_w2n_cmd_lock                 ),
  .o_icb_cmd_excl                 (slv_grp3_p0_w2n_cmd_excl                 ),
  .o_icb_cmd_xlen                 (slv_grp3_p0_w2n_cmd_xlen      [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp3_p0_w2n_cmd_xburst    [   1:   0]),
  .o_icb_cmd_modes                (slv_grp3_p0_w2n_cmd_modes     [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp3_p0_w2n_cmd_dmode                ),
  .o_icb_cmd_attri                (slv_grp3_p0_w2n_cmd_attri     [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp3_p0_w2n_cmd_beat      [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp3_p0_w2n_cmd_usr       [   2:   0]),
  .o_icb_rsp_ready                (slv_grp3_p0_w2n_rsp_ready                ),
  .o_icb_rsp_valid                (slv_grp3_p0_w2n_rsp_valid                ),
  .o_icb_rsp_err                  (slv_grp3_p0_w2n_rsp_err                  ),
  .o_icb_rsp_excl_ok              (slv_grp3_p0_w2n_rsp_excl_ok              ),
  .o_icb_rsp_rdata                (slv_grp3_p0_w2n_rsp_rdata     [  31:   0]),
  .o_icb_rsp_usr                  (slv_grp3_p0_w2n_rsp_usr       [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      assign slv_grp3_p0_w2n_rsp_usr = 3'b0;
      wire qspi0_ro_icb_bus_pend_active = 1'b0;
      wire qspi0_ro_icb_bus_icb_active;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(5+1)
      )u_qspi0_ro_icb__icb_active (
         .icb_active(qspi0_ro_icb_bus_icb_active),
            .icb_cmd_valid(slv_grp3_p0_w2n_cmd_valid),
            .icb_cmd_ready(slv_grp3_p0_w2n_cmd_ready),
            .icb_rsp_valid(slv_grp3_p0_w2n_rsp_valid),
            .icb_rsp_ready(slv_grp3_p0_w2n_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] qspi0_ro_icb_cmd_addr_full;
      assign qspi0_ro_icb_cmd_addr = qspi0_ro_icb_cmd_addr_full[32-1:0];
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(0),
    .O_SUPPORT_RATIO(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
    .OUTS_CNT_W   (5),
    .AW    (32),
    .DW    (32),
            .CMD_DP    (1),
            .RSP_DP    (1),
            .RSP_BYPBUF(0),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(1),
    .CMD_UW (1),
    .RSP_UW (1)
  )u_qspi0_ro_icb_icb_buffer(
    .i_clk_en (1'b1),
    .o_clk_en (1'b1),
    .icb_buffer_active   (),
             .i_icb_cmd_usr(1'b0),
             .i_icb_rsp_usr(),
      .i_icb_cmd_valid                (slv_grp3_p0_w2n_cmd_valid                ),
  .i_icb_cmd_ready                (slv_grp3_p0_w2n_cmd_ready                ),
  .i_icb_cmd_sel                  (slv_grp3_p0_w2n_cmd_sel                  ),
  .i_icb_cmd_read                 (slv_grp3_p0_w2n_cmd_read                 ),
  .i_icb_cmd_addr                 (slv_grp3_p0_w2n_cmd_addr      [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp3_p0_w2n_cmd_wdata     [  31:   0]),
  .i_icb_cmd_wmask                (slv_grp3_p0_w2n_cmd_wmask     [   3:   0]),
  .i_icb_cmd_size                 (slv_grp3_p0_w2n_cmd_size      [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp3_p0_w2n_cmd_lock                 ),
  .i_icb_cmd_excl                 (slv_grp3_p0_w2n_cmd_excl                 ),
  .i_icb_cmd_xlen                 (slv_grp3_p0_w2n_cmd_xlen      [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp3_p0_w2n_cmd_xburst    [   1:   0]),
  .i_icb_cmd_modes                (slv_grp3_p0_w2n_cmd_modes     [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp3_p0_w2n_cmd_dmode                ),
  .i_icb_cmd_attri                (slv_grp3_p0_w2n_cmd_attri     [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp3_p0_w2n_cmd_beat      [   1:   0]),
  .i_icb_rsp_ready                (slv_grp3_p0_w2n_rsp_ready                ),
  .i_icb_rsp_valid                (slv_grp3_p0_w2n_rsp_valid                ),
  .i_icb_rsp_err                  (slv_grp3_p0_w2n_rsp_err                  ),
  .i_icb_rsp_excl_ok              (slv_grp3_p0_w2n_rsp_excl_ok              ),
  .i_icb_rsp_rdata                (slv_grp3_p0_w2n_rsp_rdata     [  31:   0]),
      .o_icb_cmd_valid                (qspi0_ro_icb_cmd_valid                   ),
  .o_icb_cmd_ready                (qspi0_ro_icb_cmd_ready                   ),
  .o_icb_cmd_sel                  (qspi0_ro_icb_cmd_sel                     ),
  .o_icb_cmd_read                 (qspi0_ro_icb_cmd_read                    ),
  .o_icb_cmd_wdata                (qspi0_ro_icb_cmd_wdata        [  31:   0]),
  .o_icb_cmd_wmask                (qspi0_ro_icb_cmd_wmask        [   3:   0]),
  .o_icb_cmd_size                 (qspi0_ro_icb_cmd_size         [   2:   0]),
  .o_icb_cmd_lock                 (qspi0_ro_icb_cmd_lock                    ),
  .o_icb_cmd_excl                 (qspi0_ro_icb_cmd_excl                    ),
  .o_icb_cmd_xlen                 (qspi0_ro_icb_cmd_xlen         [   7:   0]),
  .o_icb_cmd_xburst               (qspi0_ro_icb_cmd_xburst       [   1:   0]),
  .o_icb_cmd_modes                (qspi0_ro_icb_cmd_modes        [   1:   0]),
  .o_icb_cmd_dmode                (qspi0_ro_icb_cmd_dmode                   ),
  .o_icb_cmd_attri                (qspi0_ro_icb_cmd_attri        [   2:   0]),
  .o_icb_cmd_beat                 (qspi0_ro_icb_cmd_beat         [   1:   0]),
  .o_icb_rsp_ready                (qspi0_ro_icb_rsp_ready                   ),
  .o_icb_rsp_valid                (qspi0_ro_icb_rsp_valid                   ),
  .o_icb_rsp_err                  (qspi0_ro_icb_rsp_err                     ),
  .o_icb_rsp_excl_ok              (qspi0_ro_icb_rsp_excl_ok                 ),
  .o_icb_rsp_rdata                (qspi0_ro_icb_rsp_rdata        [  31:   0]),
            .o_icb_cmd_usr(),
            .o_icb_rsp_usr(1'b0),
      .o_icb_cmd_addr(qspi0_ro_icb_cmd_addr_full),
      .clk  (clk_fab),  
      .rst_n(rst_n)
  );
      wire                slv_grp_4_icb_cmd_valid       ;
  wire                slv_grp_4_icb_cmd_ready       ;
  wire                slv_grp_4_icb_cmd_sel         ;
  wire                slv_grp_4_icb_cmd_read        ;
  wire    [  31:   0] slv_grp_4_icb_cmd_addr        ;
  wire    [  63:   0] slv_grp_4_icb_cmd_wdata       ;
  wire    [   7:   0] slv_grp_4_icb_cmd_wmask       ;
  wire    [   2:   0] slv_grp_4_icb_cmd_size        ;
  wire                slv_grp_4_icb_cmd_lock        ;
  wire                slv_grp_4_icb_cmd_excl        ;
  wire    [   7:   0] slv_grp_4_icb_cmd_xlen        ;
  wire    [   1:   0] slv_grp_4_icb_cmd_xburst      ;
  wire    [   1:   0] slv_grp_4_icb_cmd_modes       ;
  wire                slv_grp_4_icb_cmd_dmode       ;
  wire    [   2:   0] slv_grp_4_icb_cmd_attri       ;
  wire    [   1:   0] slv_grp_4_icb_cmd_beat        ;
  wire    [   2:   0] slv_grp_4_icb_cmd_usr         ;
  wire                slv_grp_4_icb_rsp_ready       ;
  wire                slv_grp_4_icb_rsp_valid       ;
  wire                slv_grp_4_icb_rsp_err         ;
  wire                slv_grp_4_icb_rsp_excl_ok     ;
  wire    [  63:   0] slv_grp_4_icb_rsp_rdata       ;
  wire    [   2:   0] slv_grp_4_icb_rsp_usr         ;
      wire                slv_grp_4_ro_icb_cmd_valid    ;
  wire                slv_grp_4_ro_icb_cmd_ready    ;
  wire                slv_grp_4_ro_icb_cmd_sel      ;
  wire                slv_grp_4_ro_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_4_ro_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_4_ro_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_4_ro_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_4_ro_icb_cmd_size     ;
  wire                slv_grp_4_ro_icb_cmd_lock     ;
  wire                slv_grp_4_ro_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_4_ro_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_4_ro_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_4_ro_icb_cmd_modes    ;
  wire                slv_grp_4_ro_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_4_ro_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_4_ro_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_4_ro_icb_cmd_usr      ;
  wire                slv_grp_4_ro_icb_rsp_ready    ;
  wire                slv_grp_4_ro_icb_rsp_valid    ;
  wire                slv_grp_4_ro_icb_rsp_err      ;
  wire                slv_grp_4_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_4_ro_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_4_ro_icb_rsp_usr      ;
      wire                slv_grp_4_wo_icb_cmd_valid    ;
  wire                slv_grp_4_wo_icb_cmd_ready    ;
  wire                slv_grp_4_wo_icb_cmd_sel      ;
  wire                slv_grp_4_wo_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_4_wo_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_4_wo_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_4_wo_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_4_wo_icb_cmd_size     ;
  wire                slv_grp_4_wo_icb_cmd_lock     ;
  wire                slv_grp_4_wo_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_4_wo_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_4_wo_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_4_wo_icb_cmd_modes    ;
  wire                slv_grp_4_wo_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_4_wo_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_4_wo_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_4_wo_icb_cmd_usr      ;
  wire                slv_grp_4_wo_icb_rsp_ready    ;
  wire                slv_grp_4_wo_icb_rsp_valid    ;
  wire                slv_grp_4_wo_icb_rsp_err      ;
  wire                slv_grp_4_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_4_wo_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_4_wo_icb_rsp_usr      ;
      wire                slv_grp4_p0_cmd_valid         ;
  wire                slv_grp4_p0_cmd_ready         ;
  wire                slv_grp4_p0_cmd_sel           ;
  wire                slv_grp4_p0_cmd_read          ;
  wire    [  31:   0] slv_grp4_p0_cmd_addr          ;
  wire    [  63:   0] slv_grp4_p0_cmd_wdata         ;
  wire    [   7:   0] slv_grp4_p0_cmd_wmask         ;
  wire    [   2:   0] slv_grp4_p0_cmd_size          ;
  wire                slv_grp4_p0_cmd_lock          ;
  wire                slv_grp4_p0_cmd_excl          ;
  wire    [   7:   0] slv_grp4_p0_cmd_xlen          ;
  wire    [   1:   0] slv_grp4_p0_cmd_xburst        ;
  wire    [   1:   0] slv_grp4_p0_cmd_modes         ;
  wire                slv_grp4_p0_cmd_dmode         ;
  wire    [   2:   0] slv_grp4_p0_cmd_attri         ;
  wire    [   1:   0] slv_grp4_p0_cmd_beat          ;
  wire    [   2:   0] slv_grp4_p0_cmd_usr           ;
  wire                slv_grp4_p0_rsp_ready         ;
  wire                slv_grp4_p0_rsp_valid         ;
  wire                slv_grp4_p0_rsp_err           ;
  wire                slv_grp4_p0_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp4_p0_rsp_rdata         ;
  wire    [   2:   0] slv_grp4_p0_rsp_usr           ;
      wire                slv_grp4_p0_w2n_cmd_valid     ;
  wire                slv_grp4_p0_w2n_cmd_ready     ;
  wire                slv_grp4_p0_w2n_cmd_sel       ;
  wire                slv_grp4_p0_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp4_p0_w2n_cmd_addr      ;
  wire    [  31:   0] slv_grp4_p0_w2n_cmd_wdata     ;
  wire    [   3:   0] slv_grp4_p0_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp4_p0_w2n_cmd_size      ;
  wire                slv_grp4_p0_w2n_cmd_lock      ;
  wire                slv_grp4_p0_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp4_p0_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp4_p0_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp4_p0_w2n_cmd_modes     ;
  wire                slv_grp4_p0_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp4_p0_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp4_p0_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp4_p0_w2n_cmd_usr       ;
  wire                slv_grp4_p0_w2n_rsp_ready     ;
  wire                slv_grp4_p0_w2n_rsp_valid     ;
  wire                slv_grp4_p0_w2n_rsp_err       ;
  wire                slv_grp4_p0_w2n_rsp_excl_ok   ;
  wire    [  31:   0] slv_grp4_p0_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp4_p0_w2n_rsp_usr       ;
      wire                slv_grp4_p0_ro_cmd_valid      ;
  wire                slv_grp4_p0_ro_cmd_ready      ;
  wire                slv_grp4_p0_ro_cmd_sel        ;
  wire                slv_grp4_p0_ro_cmd_read       ;
  wire    [  31:   0] slv_grp4_p0_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp4_p0_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp4_p0_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp4_p0_ro_cmd_size       ;
  wire                slv_grp4_p0_ro_cmd_lock       ;
  wire                slv_grp4_p0_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp4_p0_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp4_p0_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp4_p0_ro_cmd_modes      ;
  wire                slv_grp4_p0_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp4_p0_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp4_p0_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp4_p0_ro_cmd_usr        ;
  wire                slv_grp4_p0_ro_rsp_ready      ;
  wire                slv_grp4_p0_ro_rsp_valid      ;
  wire                slv_grp4_p0_ro_rsp_err        ;
  wire                slv_grp4_p0_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp4_p0_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp4_p0_ro_rsp_usr        ;
      wire                slv_grp4_p0_w2n_ro_cmd_valid  ;
  wire                slv_grp4_p0_w2n_ro_cmd_ready  ;
  wire                slv_grp4_p0_w2n_ro_cmd_sel    ;
  wire                slv_grp4_p0_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp4_p0_w2n_ro_cmd_addr   ;
  wire    [  31:   0] slv_grp4_p0_w2n_ro_cmd_wdata  ;
  wire    [   3:   0] slv_grp4_p0_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp4_p0_w2n_ro_cmd_size   ;
  wire                slv_grp4_p0_w2n_ro_cmd_lock   ;
  wire                slv_grp4_p0_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp4_p0_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp4_p0_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp4_p0_w2n_ro_cmd_modes  ;
  wire                slv_grp4_p0_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp4_p0_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp4_p0_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp4_p0_w2n_ro_cmd_usr    ;
  wire                slv_grp4_p0_w2n_ro_rsp_ready  ;
  wire                slv_grp4_p0_w2n_ro_rsp_valid  ;
  wire                slv_grp4_p0_w2n_ro_rsp_err    ;
  wire                slv_grp4_p0_w2n_ro_rsp_excl_ok ;
  wire    [  31:   0] slv_grp4_p0_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp4_p0_w2n_ro_rsp_usr    ;
      wire                slv_grp4_p0_wo_cmd_valid      ;
  wire                slv_grp4_p0_wo_cmd_ready      ;
  wire                slv_grp4_p0_wo_cmd_sel        ;
  wire                slv_grp4_p0_wo_cmd_read       ;
  wire    [  31:   0] slv_grp4_p0_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp4_p0_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp4_p0_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp4_p0_wo_cmd_size       ;
  wire                slv_grp4_p0_wo_cmd_lock       ;
  wire                slv_grp4_p0_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp4_p0_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp4_p0_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp4_p0_wo_cmd_modes      ;
  wire                slv_grp4_p0_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp4_p0_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp4_p0_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp4_p0_wo_cmd_usr        ;
  wire                slv_grp4_p0_wo_rsp_ready      ;
  wire                slv_grp4_p0_wo_rsp_valid      ;
  wire                slv_grp4_p0_wo_rsp_err        ;
  wire                slv_grp4_p0_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp4_p0_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp4_p0_wo_rsp_usr        ;
      wire                slv_grp4_p0_w2n_wo_cmd_valid  ;
  wire                slv_grp4_p0_w2n_wo_cmd_ready  ;
  wire                slv_grp4_p0_w2n_wo_cmd_sel    ;
  wire                slv_grp4_p0_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp4_p0_w2n_wo_cmd_addr   ;
  wire    [  31:   0] slv_grp4_p0_w2n_wo_cmd_wdata  ;
  wire    [   3:   0] slv_grp4_p0_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp4_p0_w2n_wo_cmd_size   ;
  wire                slv_grp4_p0_w2n_wo_cmd_lock   ;
  wire                slv_grp4_p0_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp4_p0_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp4_p0_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp4_p0_w2n_wo_cmd_modes  ;
  wire                slv_grp4_p0_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp4_p0_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp4_p0_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp4_p0_w2n_wo_cmd_usr    ;
  wire                slv_grp4_p0_w2n_wo_rsp_ready  ;
  wire                slv_grp4_p0_w2n_wo_rsp_valid  ;
  wire                slv_grp4_p0_w2n_wo_rsp_err    ;
  wire                slv_grp4_p0_w2n_wo_rsp_excl_ok ;
  wire    [  31:   0] slv_grp4_p0_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp4_p0_w2n_wo_rsp_usr    ;
                wire                      slv_grp4_p0_w2n_wo_rsp_last;
      wire                slv_grp4_p1_cmd_valid         ;
  wire                slv_grp4_p1_cmd_ready         ;
  wire                slv_grp4_p1_cmd_sel           ;
  wire                slv_grp4_p1_cmd_read          ;
  wire    [  31:   0] slv_grp4_p1_cmd_addr          ;
  wire    [  63:   0] slv_grp4_p1_cmd_wdata         ;
  wire    [   7:   0] slv_grp4_p1_cmd_wmask         ;
  wire    [   2:   0] slv_grp4_p1_cmd_size          ;
  wire                slv_grp4_p1_cmd_lock          ;
  wire                slv_grp4_p1_cmd_excl          ;
  wire    [   7:   0] slv_grp4_p1_cmd_xlen          ;
  wire    [   1:   0] slv_grp4_p1_cmd_xburst        ;
  wire    [   1:   0] slv_grp4_p1_cmd_modes         ;
  wire                slv_grp4_p1_cmd_dmode         ;
  wire    [   2:   0] slv_grp4_p1_cmd_attri         ;
  wire    [   1:   0] slv_grp4_p1_cmd_beat          ;
  wire    [   2:   0] slv_grp4_p1_cmd_usr           ;
  wire                slv_grp4_p1_rsp_ready         ;
  wire                slv_grp4_p1_rsp_valid         ;
  wire                slv_grp4_p1_rsp_err           ;
  wire                slv_grp4_p1_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp4_p1_rsp_rdata         ;
  wire    [   2:   0] slv_grp4_p1_rsp_usr           ;
      wire                slv_grp4_p1_w2n_cmd_valid     ;
  wire                slv_grp4_p1_w2n_cmd_ready     ;
  wire                slv_grp4_p1_w2n_cmd_sel       ;
  wire                slv_grp4_p1_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp4_p1_w2n_cmd_addr      ;
  wire    [  31:   0] slv_grp4_p1_w2n_cmd_wdata     ;
  wire    [   3:   0] slv_grp4_p1_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp4_p1_w2n_cmd_size      ;
  wire                slv_grp4_p1_w2n_cmd_lock      ;
  wire                slv_grp4_p1_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp4_p1_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp4_p1_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp4_p1_w2n_cmd_modes     ;
  wire                slv_grp4_p1_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp4_p1_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp4_p1_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp4_p1_w2n_cmd_usr       ;
  wire                slv_grp4_p1_w2n_rsp_ready     ;
  wire                slv_grp4_p1_w2n_rsp_valid     ;
  wire                slv_grp4_p1_w2n_rsp_err       ;
  wire                slv_grp4_p1_w2n_rsp_excl_ok   ;
  wire    [  31:   0] slv_grp4_p1_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp4_p1_w2n_rsp_usr       ;
      wire                slv_grp4_p1_ro_cmd_valid      ;
  wire                slv_grp4_p1_ro_cmd_ready      ;
  wire                slv_grp4_p1_ro_cmd_sel        ;
  wire                slv_grp4_p1_ro_cmd_read       ;
  wire    [  31:   0] slv_grp4_p1_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp4_p1_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp4_p1_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp4_p1_ro_cmd_size       ;
  wire                slv_grp4_p1_ro_cmd_lock       ;
  wire                slv_grp4_p1_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp4_p1_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp4_p1_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp4_p1_ro_cmd_modes      ;
  wire                slv_grp4_p1_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp4_p1_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp4_p1_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp4_p1_ro_cmd_usr        ;
  wire                slv_grp4_p1_ro_rsp_ready      ;
  wire                slv_grp4_p1_ro_rsp_valid      ;
  wire                slv_grp4_p1_ro_rsp_err        ;
  wire                slv_grp4_p1_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp4_p1_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp4_p1_ro_rsp_usr        ;
      wire                slv_grp4_p1_w2n_ro_cmd_valid  ;
  wire                slv_grp4_p1_w2n_ro_cmd_ready  ;
  wire                slv_grp4_p1_w2n_ro_cmd_sel    ;
  wire                slv_grp4_p1_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp4_p1_w2n_ro_cmd_addr   ;
  wire    [  31:   0] slv_grp4_p1_w2n_ro_cmd_wdata  ;
  wire    [   3:   0] slv_grp4_p1_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp4_p1_w2n_ro_cmd_size   ;
  wire                slv_grp4_p1_w2n_ro_cmd_lock   ;
  wire                slv_grp4_p1_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp4_p1_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp4_p1_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp4_p1_w2n_ro_cmd_modes  ;
  wire                slv_grp4_p1_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp4_p1_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp4_p1_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp4_p1_w2n_ro_cmd_usr    ;
  wire                slv_grp4_p1_w2n_ro_rsp_ready  ;
  wire                slv_grp4_p1_w2n_ro_rsp_valid  ;
  wire                slv_grp4_p1_w2n_ro_rsp_err    ;
  wire                slv_grp4_p1_w2n_ro_rsp_excl_ok ;
  wire    [  31:   0] slv_grp4_p1_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp4_p1_w2n_ro_rsp_usr    ;
      wire                slv_grp4_p1_wo_cmd_valid      ;
  wire                slv_grp4_p1_wo_cmd_ready      ;
  wire                slv_grp4_p1_wo_cmd_sel        ;
  wire                slv_grp4_p1_wo_cmd_read       ;
  wire    [  31:   0] slv_grp4_p1_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp4_p1_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp4_p1_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp4_p1_wo_cmd_size       ;
  wire                slv_grp4_p1_wo_cmd_lock       ;
  wire                slv_grp4_p1_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp4_p1_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp4_p1_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp4_p1_wo_cmd_modes      ;
  wire                slv_grp4_p1_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp4_p1_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp4_p1_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp4_p1_wo_cmd_usr        ;
  wire                slv_grp4_p1_wo_rsp_ready      ;
  wire                slv_grp4_p1_wo_rsp_valid      ;
  wire                slv_grp4_p1_wo_rsp_err        ;
  wire                slv_grp4_p1_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp4_p1_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp4_p1_wo_rsp_usr        ;
      wire                slv_grp4_p1_w2n_wo_cmd_valid  ;
  wire                slv_grp4_p1_w2n_wo_cmd_ready  ;
  wire                slv_grp4_p1_w2n_wo_cmd_sel    ;
  wire                slv_grp4_p1_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp4_p1_w2n_wo_cmd_addr   ;
  wire    [  31:   0] slv_grp4_p1_w2n_wo_cmd_wdata  ;
  wire    [   3:   0] slv_grp4_p1_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp4_p1_w2n_wo_cmd_size   ;
  wire                slv_grp4_p1_w2n_wo_cmd_lock   ;
  wire                slv_grp4_p1_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp4_p1_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp4_p1_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp4_p1_w2n_wo_cmd_modes  ;
  wire                slv_grp4_p1_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp4_p1_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp4_p1_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp4_p1_w2n_wo_cmd_usr    ;
  wire                slv_grp4_p1_w2n_wo_rsp_ready  ;
  wire                slv_grp4_p1_w2n_wo_rsp_valid  ;
  wire                slv_grp4_p1_w2n_wo_rsp_err    ;
  wire                slv_grp4_p1_w2n_wo_rsp_excl_ok ;
  wire    [  31:   0] slv_grp4_p1_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp4_p1_w2n_wo_rsp_usr    ;
                wire                      slv_grp4_p1_w2n_wo_rsp_last;
   e603_subsys_sgrp4_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (32'h10000000 + 32'h2000),
      .O0_BASE_REGION_LSB(12),
      .O1_BASE_ADDR      (32'h10000000),
      .O1_BASE_REGION_LSB(20),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (16 ),
      .SPLT_FIFO_OUTS_CNT_W(5),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp4_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_4_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (slv_grp_4_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (slv_grp_4_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (slv_grp_4_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (slv_grp_4_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_4_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_4_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_4_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_4_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (slv_grp_4_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (slv_grp_4_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_4_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_4_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_4_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (slv_grp_4_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_4_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_4_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_4_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (slv_grp_4_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (slv_grp_4_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (slv_grp_4_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (slv_grp_4_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_4_icb_rsp_usr         [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (slv_grp4_p0_cmd_valid                    ),
  .o0_icb_cmd_ready               (slv_grp4_p0_cmd_ready                    ),
  .o0_icb_cmd_sel                 (slv_grp4_p0_cmd_sel                      ),
  .o0_icb_cmd_read                (slv_grp4_p0_cmd_read                     ),
  .o0_icb_cmd_addr                (slv_grp4_p0_cmd_addr          [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp4_p0_cmd_wdata         [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp4_p0_cmd_wmask         [   7:   0]),
  .o0_icb_cmd_size                (slv_grp4_p0_cmd_size          [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp4_p0_cmd_lock                     ),
  .o0_icb_cmd_excl                (slv_grp4_p0_cmd_excl                     ),
  .o0_icb_cmd_xlen                (slv_grp4_p0_cmd_xlen          [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp4_p0_cmd_xburst        [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp4_p0_cmd_modes         [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp4_p0_cmd_dmode                    ),
  .o0_icb_cmd_attri               (slv_grp4_p0_cmd_attri         [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp4_p0_cmd_beat          [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp4_p0_cmd_usr           [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp4_p0_rsp_ready                    ),
  .o0_icb_rsp_valid               (slv_grp4_p0_rsp_valid                    ),
  .o0_icb_rsp_err                 (slv_grp4_p0_rsp_err                      ),
  .o0_icb_rsp_excl_ok             (slv_grp4_p0_rsp_excl_ok                  ),
  .o0_icb_rsp_rdata               (slv_grp4_p0_rsp_rdata         [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp4_p0_rsp_usr           [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (slv_grp4_p1_cmd_valid                    ),
  .o1_icb_cmd_ready               (slv_grp4_p1_cmd_ready                    ),
  .o1_icb_cmd_sel                 (slv_grp4_p1_cmd_sel                      ),
  .o1_icb_cmd_read                (slv_grp4_p1_cmd_read                     ),
  .o1_icb_cmd_addr                (slv_grp4_p1_cmd_addr          [  31:   0]),
  .o1_icb_cmd_wdata               (slv_grp4_p1_cmd_wdata         [  63:   0]),
  .o1_icb_cmd_wmask               (slv_grp4_p1_cmd_wmask         [   7:   0]),
  .o1_icb_cmd_size                (slv_grp4_p1_cmd_size          [   2:   0]),
  .o1_icb_cmd_lock                (slv_grp4_p1_cmd_lock                     ),
  .o1_icb_cmd_excl                (slv_grp4_p1_cmd_excl                     ),
  .o1_icb_cmd_xlen                (slv_grp4_p1_cmd_xlen          [   7:   0]),
  .o1_icb_cmd_xburst              (slv_grp4_p1_cmd_xburst        [   1:   0]),
  .o1_icb_cmd_modes               (slv_grp4_p1_cmd_modes         [   1:   0]),
  .o1_icb_cmd_dmode               (slv_grp4_p1_cmd_dmode                    ),
  .o1_icb_cmd_attri               (slv_grp4_p1_cmd_attri         [   2:   0]),
  .o1_icb_cmd_beat                (slv_grp4_p1_cmd_beat          [   1:   0]),
  .o1_icb_cmd_usr                 (slv_grp4_p1_cmd_usr           [   2:   0]),
  .o1_icb_rsp_ready               (slv_grp4_p1_rsp_ready                    ),
  .o1_icb_rsp_valid               (slv_grp4_p1_rsp_valid                    ),
  .o1_icb_rsp_err                 (slv_grp4_p1_rsp_err                      ),
  .o1_icb_rsp_excl_ok             (slv_grp4_p1_rsp_excl_ok                  ),
  .o1_icb_rsp_rdata               (slv_grp4_p1_rsp_rdata         [  63:   0]),
  .o1_icb_rsp_usr                 (slv_grp4_p1_rsp_usr           [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (16),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(32 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_eth_cfg_apb_icb_wconv(
        .i_icb_cmd_valid                (slv_grp4_p0_cmd_valid                    ),
  .i_icb_cmd_ready                (slv_grp4_p0_cmd_ready                    ),
  .i_icb_cmd_sel                  (slv_grp4_p0_cmd_sel                      ),
  .i_icb_cmd_read                 (slv_grp4_p0_cmd_read                     ),
  .i_icb_cmd_addr                 (slv_grp4_p0_cmd_addr          [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp4_p0_cmd_wdata         [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp4_p0_cmd_wmask         [   7:   0]),
  .i_icb_cmd_size                 (slv_grp4_p0_cmd_size          [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp4_p0_cmd_lock                     ),
  .i_icb_cmd_excl                 (slv_grp4_p0_cmd_excl                     ),
  .i_icb_cmd_xlen                 (slv_grp4_p0_cmd_xlen          [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp4_p0_cmd_xburst        [   1:   0]),
  .i_icb_cmd_modes                (slv_grp4_p0_cmd_modes         [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp4_p0_cmd_dmode                    ),
  .i_icb_cmd_attri                (slv_grp4_p0_cmd_attri         [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp4_p0_cmd_beat          [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp4_p0_cmd_usr           [   2:   0]),
  .i_icb_rsp_ready                (slv_grp4_p0_rsp_ready                    ),
  .i_icb_rsp_valid                (slv_grp4_p0_rsp_valid                    ),
  .i_icb_rsp_err                  (slv_grp4_p0_rsp_err                      ),
  .i_icb_rsp_excl_ok              (slv_grp4_p0_rsp_excl_ok                  ),
  .i_icb_rsp_rdata                (slv_grp4_p0_rsp_rdata         [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp4_p0_rsp_usr           [   2:   0]),
        .o_icb_cmd_valid                (slv_grp4_p0_w2n_cmd_valid                ),
  .o_icb_cmd_ready                (slv_grp4_p0_w2n_cmd_ready                ),
  .o_icb_cmd_sel                  (slv_grp4_p0_w2n_cmd_sel                  ),
  .o_icb_cmd_read                 (slv_grp4_p0_w2n_cmd_read                 ),
  .o_icb_cmd_addr                 (slv_grp4_p0_w2n_cmd_addr      [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp4_p0_w2n_cmd_wdata     [  31:   0]),
  .o_icb_cmd_wmask                (slv_grp4_p0_w2n_cmd_wmask     [   3:   0]),
  .o_icb_cmd_size                 (slv_grp4_p0_w2n_cmd_size      [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp4_p0_w2n_cmd_lock                 ),
  .o_icb_cmd_excl                 (slv_grp4_p0_w2n_cmd_excl                 ),
  .o_icb_cmd_xlen                 (slv_grp4_p0_w2n_cmd_xlen      [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp4_p0_w2n_cmd_xburst    [   1:   0]),
  .o_icb_cmd_modes                (slv_grp4_p0_w2n_cmd_modes     [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp4_p0_w2n_cmd_dmode                ),
  .o_icb_cmd_attri                (slv_grp4_p0_w2n_cmd_attri     [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp4_p0_w2n_cmd_beat      [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp4_p0_w2n_cmd_usr       [   2:   0]),
  .o_icb_rsp_ready                (slv_grp4_p0_w2n_rsp_ready                ),
  .o_icb_rsp_valid                (slv_grp4_p0_w2n_rsp_valid                ),
  .o_icb_rsp_err                  (slv_grp4_p0_w2n_rsp_err                  ),
  .o_icb_rsp_excl_ok              (slv_grp4_p0_w2n_rsp_excl_ok              ),
  .o_icb_rsp_rdata                (slv_grp4_p0_w2n_rsp_rdata     [  31:   0]),
  .o_icb_rsp_usr                  (slv_grp4_p0_w2n_rsp_usr       [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      wire eth_cfg_apb_bus_pend_active = 1'b0;
            wire eth_cfg_apb_bus_icb_active;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(5+1)
      )u_eth_cfg_apb__icb_active (
         .icb_active(eth_cfg_apb_bus_icb_active),
            .icb_cmd_valid(slv_grp4_p0_w2n_cmd_valid),
            .icb_cmd_ready(slv_grp4_p0_w2n_cmd_ready),
            .icb_rsp_valid(slv_grp4_p0_w2n_rsp_valid),
            .icb_rsp_ready(slv_grp4_p0_w2n_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire[32-1:0] eth_cfg_apb_paddr_full;
      assign eth_cfg_apb_paddr = eth_cfg_apb_paddr_full[12-1:0];
      assign slv_grp4_p0_w2n_rsp_usr = 3'b0;
  e603_subsys_gnrl_usr_ficb2apb_ratio # (
    .OUTS_CNT_W(5),
      .SUPPORT_RATIO(0), 
      .CMD_DP    (1),
      .RSP_DP    (1),
      .RSP_BYPBUF(0),
      .AW(32),
      .DW(32) 
    ) u_eth_cfg_apb_icb2apb_ratio(
    .ratio_apb_clk_en (1'b1),
    .icb_clk_en (1'b1),
    .icb2apb_ratio_active(),
      .icb_cmd_valid                  (slv_grp4_p0_w2n_cmd_valid                ),
  .icb_cmd_ready                  (slv_grp4_p0_w2n_cmd_ready                ),
  .icb_cmd_sel                    (slv_grp4_p0_w2n_cmd_sel                  ),
  .icb_cmd_read                   (slv_grp4_p0_w2n_cmd_read                 ),
  .icb_cmd_wdata                  (slv_grp4_p0_w2n_cmd_wdata     [  31:   0]),
  .icb_cmd_wmask                  (slv_grp4_p0_w2n_cmd_wmask     [   3:   0]),
  .icb_cmd_size                   (slv_grp4_p0_w2n_cmd_size      [   2:   0]),
  .icb_cmd_lock                   (slv_grp4_p0_w2n_cmd_lock                 ),
  .icb_cmd_excl                   (slv_grp4_p0_w2n_cmd_excl                 ),
  .icb_cmd_xlen                   (slv_grp4_p0_w2n_cmd_xlen      [   7:   0]),
  .icb_cmd_xburst                 (slv_grp4_p0_w2n_cmd_xburst    [   1:   0]),
  .icb_cmd_modes                  (slv_grp4_p0_w2n_cmd_modes     [   1:   0]),
  .icb_cmd_dmode                  (slv_grp4_p0_w2n_cmd_dmode                ),
  .icb_cmd_attri                  (slv_grp4_p0_w2n_cmd_attri     [   2:   0]),
  .icb_cmd_beat                   (slv_grp4_p0_w2n_cmd_beat      [   1:   0]),
  .icb_rsp_ready                  (slv_grp4_p0_w2n_rsp_ready                ),
  .icb_rsp_valid                  (slv_grp4_p0_w2n_rsp_valid                ),
  .icb_rsp_err                    (slv_grp4_p0_w2n_rsp_err                  ),
  .icb_rsp_excl_ok                (slv_grp4_p0_w2n_rsp_excl_ok              ),
  .icb_rsp_rdata                  (slv_grp4_p0_w2n_rsp_rdata     [  31:   0]),
      .icb_cmd_addr(slv_grp4_p0_w2n_cmd_addr),
      .ratio_apb_pwrite               (eth_cfg_apb_pwrite                       ),
  .ratio_apb_psel                 (eth_cfg_apb_psel                         ),
  .ratio_apb_pprot                (eth_cfg_apb_pprot             [   2:   0]),
  .ratio_apb_pstrobe              (eth_cfg_apb_pstrobe           [   3:   0]),
  .ratio_apb_penable              (eth_cfg_apb_penable                      ),
  .ratio_apb_pwdata               (eth_cfg_apb_pwdata            [  31:   0]),
  .ratio_apb_prdata               (eth_cfg_apb_prdata            [  31:   0]),
  .ratio_apb_pready               (eth_cfg_apb_pready                       ),
  .ratio_apb_pslverr              (eth_cfg_apb_pslverr                      ),
      .ratio_apb_paddr(eth_cfg_apb_paddr_full),
      .icb_cmd_usr(1'b0),
      .icb_rsp_usr(),
            .ratio_apb_puser (),
            .ratio_apb_pruser(1'b0),
    .clk            (clk_fab  ),
    .rst_n          (rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (16),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(32 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_biu2ppi_icb_icb_wconv(
        .i_icb_cmd_valid                (slv_grp4_p1_cmd_valid                    ),
  .i_icb_cmd_ready                (slv_grp4_p1_cmd_ready                    ),
  .i_icb_cmd_sel                  (slv_grp4_p1_cmd_sel                      ),
  .i_icb_cmd_read                 (slv_grp4_p1_cmd_read                     ),
  .i_icb_cmd_addr                 (slv_grp4_p1_cmd_addr          [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp4_p1_cmd_wdata         [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp4_p1_cmd_wmask         [   7:   0]),
  .i_icb_cmd_size                 (slv_grp4_p1_cmd_size          [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp4_p1_cmd_lock                     ),
  .i_icb_cmd_excl                 (slv_grp4_p1_cmd_excl                     ),
  .i_icb_cmd_xlen                 (slv_grp4_p1_cmd_xlen          [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp4_p1_cmd_xburst        [   1:   0]),
  .i_icb_cmd_modes                (slv_grp4_p1_cmd_modes         [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp4_p1_cmd_dmode                    ),
  .i_icb_cmd_attri                (slv_grp4_p1_cmd_attri         [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp4_p1_cmd_beat          [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp4_p1_cmd_usr           [   2:   0]),
  .i_icb_rsp_ready                (slv_grp4_p1_rsp_ready                    ),
  .i_icb_rsp_valid                (slv_grp4_p1_rsp_valid                    ),
  .i_icb_rsp_err                  (slv_grp4_p1_rsp_err                      ),
  .i_icb_rsp_excl_ok              (slv_grp4_p1_rsp_excl_ok                  ),
  .i_icb_rsp_rdata                (slv_grp4_p1_rsp_rdata         [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp4_p1_rsp_usr           [   2:   0]),
        .o_icb_cmd_valid                (slv_grp4_p1_w2n_cmd_valid                ),
  .o_icb_cmd_ready                (slv_grp4_p1_w2n_cmd_ready                ),
  .o_icb_cmd_sel                  (slv_grp4_p1_w2n_cmd_sel                  ),
  .o_icb_cmd_read                 (slv_grp4_p1_w2n_cmd_read                 ),
  .o_icb_cmd_addr                 (slv_grp4_p1_w2n_cmd_addr      [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp4_p1_w2n_cmd_wdata     [  31:   0]),
  .o_icb_cmd_wmask                (slv_grp4_p1_w2n_cmd_wmask     [   3:   0]),
  .o_icb_cmd_size                 (slv_grp4_p1_w2n_cmd_size      [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp4_p1_w2n_cmd_lock                 ),
  .o_icb_cmd_excl                 (slv_grp4_p1_w2n_cmd_excl                 ),
  .o_icb_cmd_xlen                 (slv_grp4_p1_w2n_cmd_xlen      [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp4_p1_w2n_cmd_xburst    [   1:   0]),
  .o_icb_cmd_modes                (slv_grp4_p1_w2n_cmd_modes     [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp4_p1_w2n_cmd_dmode                ),
  .o_icb_cmd_attri                (slv_grp4_p1_w2n_cmd_attri     [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp4_p1_w2n_cmd_beat      [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp4_p1_w2n_cmd_usr       [   2:   0]),
  .o_icb_rsp_ready                (slv_grp4_p1_w2n_rsp_ready                ),
  .o_icb_rsp_valid                (slv_grp4_p1_w2n_rsp_valid                ),
  .o_icb_rsp_err                  (slv_grp4_p1_w2n_rsp_err                  ),
  .o_icb_rsp_excl_ok              (slv_grp4_p1_w2n_rsp_excl_ok              ),
  .o_icb_rsp_rdata                (slv_grp4_p1_w2n_rsp_rdata     [  31:   0]),
  .o_icb_rsp_usr                  (slv_grp4_p1_w2n_rsp_usr       [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      assign slv_grp4_p1_w2n_rsp_usr = 3'b0;
      wire biu2ppi_icb_bus_pend_active = 1'b0;
      wire biu2ppi_icb_bus_icb_active;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(5+1)
      )u_biu2ppi_icb__icb_active (
         .icb_active(biu2ppi_icb_bus_icb_active),
            .icb_cmd_valid(slv_grp4_p1_w2n_cmd_valid),
            .icb_cmd_ready(slv_grp4_p1_w2n_cmd_ready),
            .icb_rsp_valid(slv_grp4_p1_w2n_rsp_valid),
            .icb_rsp_ready(slv_grp4_p1_w2n_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] biu2ppi_icb_cmd_addr_full;
      assign biu2ppi_icb_cmd_addr = biu2ppi_icb_cmd_addr_full[32-1:0];
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(0),
    .O_SUPPORT_RATIO(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
    .OUTS_CNT_W   (5),
    .AW    (32),
    .DW    (32),
            .CMD_DP    (2),
            .RSP_DP    (2),
            .RSP_BYPBUF(0),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(0),
    .CMD_UW (1),
    .RSP_UW (1)
  )u_biu2ppi_icb_icb_buffer(
    .i_clk_en (1'b1),
    .o_clk_en (1'b1),
    .icb_buffer_active   (),
             .i_icb_cmd_usr(1'b0),
             .i_icb_rsp_usr(),
      .i_icb_cmd_valid                (slv_grp4_p1_w2n_cmd_valid                ),
  .i_icb_cmd_ready                (slv_grp4_p1_w2n_cmd_ready                ),
  .i_icb_cmd_sel                  (slv_grp4_p1_w2n_cmd_sel                  ),
  .i_icb_cmd_read                 (slv_grp4_p1_w2n_cmd_read                 ),
  .i_icb_cmd_addr                 (slv_grp4_p1_w2n_cmd_addr      [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp4_p1_w2n_cmd_wdata     [  31:   0]),
  .i_icb_cmd_wmask                (slv_grp4_p1_w2n_cmd_wmask     [   3:   0]),
  .i_icb_cmd_size                 (slv_grp4_p1_w2n_cmd_size      [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp4_p1_w2n_cmd_lock                 ),
  .i_icb_cmd_excl                 (slv_grp4_p1_w2n_cmd_excl                 ),
  .i_icb_cmd_xlen                 (slv_grp4_p1_w2n_cmd_xlen      [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp4_p1_w2n_cmd_xburst    [   1:   0]),
  .i_icb_cmd_modes                (slv_grp4_p1_w2n_cmd_modes     [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp4_p1_w2n_cmd_dmode                ),
  .i_icb_cmd_attri                (slv_grp4_p1_w2n_cmd_attri     [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp4_p1_w2n_cmd_beat      [   1:   0]),
  .i_icb_rsp_ready                (slv_grp4_p1_w2n_rsp_ready                ),
  .i_icb_rsp_valid                (slv_grp4_p1_w2n_rsp_valid                ),
  .i_icb_rsp_err                  (slv_grp4_p1_w2n_rsp_err                  ),
  .i_icb_rsp_excl_ok              (slv_grp4_p1_w2n_rsp_excl_ok              ),
  .i_icb_rsp_rdata                (slv_grp4_p1_w2n_rsp_rdata     [  31:   0]),
      .o_icb_cmd_valid                (biu2ppi_icb_cmd_valid                    ),
  .o_icb_cmd_ready                (biu2ppi_icb_cmd_ready                    ),
  .o_icb_cmd_sel                  (biu2ppi_icb_cmd_sel                      ),
  .o_icb_cmd_read                 (biu2ppi_icb_cmd_read                     ),
  .o_icb_cmd_wdata                (biu2ppi_icb_cmd_wdata         [  31:   0]),
  .o_icb_cmd_wmask                (biu2ppi_icb_cmd_wmask         [   3:   0]),
  .o_icb_cmd_size                 (biu2ppi_icb_cmd_size          [   2:   0]),
  .o_icb_cmd_lock                 (biu2ppi_icb_cmd_lock                     ),
  .o_icb_cmd_excl                 (biu2ppi_icb_cmd_excl                     ),
  .o_icb_cmd_xlen                 (biu2ppi_icb_cmd_xlen          [   7:   0]),
  .o_icb_cmd_xburst               (biu2ppi_icb_cmd_xburst        [   1:   0]),
  .o_icb_cmd_modes                (biu2ppi_icb_cmd_modes         [   1:   0]),
  .o_icb_cmd_dmode                (biu2ppi_icb_cmd_dmode                    ),
  .o_icb_cmd_attri                (biu2ppi_icb_cmd_attri         [   2:   0]),
  .o_icb_cmd_beat                 (biu2ppi_icb_cmd_beat          [   1:   0]),
  .o_icb_rsp_ready                (biu2ppi_icb_rsp_ready                    ),
  .o_icb_rsp_valid                (biu2ppi_icb_rsp_valid                    ),
  .o_icb_rsp_err                  (biu2ppi_icb_rsp_err                      ),
  .o_icb_rsp_excl_ok              (biu2ppi_icb_rsp_excl_ok                  ),
  .o_icb_rsp_rdata                (biu2ppi_icb_rsp_rdata         [  31:   0]),
            .o_icb_cmd_usr(),
            .o_icb_rsp_usr(1'b0),
      .o_icb_cmd_addr(biu2ppi_icb_cmd_addr_full),
      .clk  (clk_fab),  
      .rst_n(rst_n)
  );
      wire                slv_grp_5_icb_cmd_valid       ;
  wire                slv_grp_5_icb_cmd_ready       ;
  wire                slv_grp_5_icb_cmd_sel         ;
  wire                slv_grp_5_icb_cmd_read        ;
  wire    [  31:   0] slv_grp_5_icb_cmd_addr        ;
  wire    [  63:   0] slv_grp_5_icb_cmd_wdata       ;
  wire    [   7:   0] slv_grp_5_icb_cmd_wmask       ;
  wire    [   2:   0] slv_grp_5_icb_cmd_size        ;
  wire                slv_grp_5_icb_cmd_lock        ;
  wire                slv_grp_5_icb_cmd_excl        ;
  wire    [   7:   0] slv_grp_5_icb_cmd_xlen        ;
  wire    [   1:   0] slv_grp_5_icb_cmd_xburst      ;
  wire    [   1:   0] slv_grp_5_icb_cmd_modes       ;
  wire                slv_grp_5_icb_cmd_dmode       ;
  wire    [   2:   0] slv_grp_5_icb_cmd_attri       ;
  wire    [   1:   0] slv_grp_5_icb_cmd_beat        ;
  wire    [   2:   0] slv_grp_5_icb_cmd_usr         ;
  wire                slv_grp_5_icb_rsp_ready       ;
  wire                slv_grp_5_icb_rsp_valid       ;
  wire                slv_grp_5_icb_rsp_err         ;
  wire                slv_grp_5_icb_rsp_excl_ok     ;
  wire    [  63:   0] slv_grp_5_icb_rsp_rdata       ;
  wire    [   2:   0] slv_grp_5_icb_rsp_usr         ;
      wire                slv_grp_5_ro_icb_cmd_valid    ;
  wire                slv_grp_5_ro_icb_cmd_ready    ;
  wire                slv_grp_5_ro_icb_cmd_sel      ;
  wire                slv_grp_5_ro_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_5_ro_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_5_ro_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_5_ro_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_5_ro_icb_cmd_size     ;
  wire                slv_grp_5_ro_icb_cmd_lock     ;
  wire                slv_grp_5_ro_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_5_ro_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_5_ro_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_5_ro_icb_cmd_modes    ;
  wire                slv_grp_5_ro_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_5_ro_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_5_ro_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_5_ro_icb_cmd_usr      ;
  wire                slv_grp_5_ro_icb_rsp_ready    ;
  wire                slv_grp_5_ro_icb_rsp_valid    ;
  wire                slv_grp_5_ro_icb_rsp_err      ;
  wire                slv_grp_5_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_5_ro_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_5_ro_icb_rsp_usr      ;
      wire                slv_grp_5_wo_icb_cmd_valid    ;
  wire                slv_grp_5_wo_icb_cmd_ready    ;
  wire                slv_grp_5_wo_icb_cmd_sel      ;
  wire                slv_grp_5_wo_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_5_wo_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_5_wo_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_5_wo_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_5_wo_icb_cmd_size     ;
  wire                slv_grp_5_wo_icb_cmd_lock     ;
  wire                slv_grp_5_wo_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_5_wo_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_5_wo_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_5_wo_icb_cmd_modes    ;
  wire                slv_grp_5_wo_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_5_wo_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_5_wo_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_5_wo_icb_cmd_usr      ;
  wire                slv_grp_5_wo_icb_rsp_ready    ;
  wire                slv_grp_5_wo_icb_rsp_valid    ;
  wire                slv_grp_5_wo_icb_rsp_err      ;
  wire                slv_grp_5_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_5_wo_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_5_wo_icb_rsp_usr      ;
      wire                slv_grp5_p0_cmd_valid         ;
  wire                slv_grp5_p0_cmd_ready         ;
  wire                slv_grp5_p0_cmd_sel           ;
  wire                slv_grp5_p0_cmd_read          ;
  wire    [  31:   0] slv_grp5_p0_cmd_addr          ;
  wire    [  63:   0] slv_grp5_p0_cmd_wdata         ;
  wire    [   7:   0] slv_grp5_p0_cmd_wmask         ;
  wire    [   2:   0] slv_grp5_p0_cmd_size          ;
  wire                slv_grp5_p0_cmd_lock          ;
  wire                slv_grp5_p0_cmd_excl          ;
  wire    [   7:   0] slv_grp5_p0_cmd_xlen          ;
  wire    [   1:   0] slv_grp5_p0_cmd_xburst        ;
  wire    [   1:   0] slv_grp5_p0_cmd_modes         ;
  wire                slv_grp5_p0_cmd_dmode         ;
  wire    [   2:   0] slv_grp5_p0_cmd_attri         ;
  wire    [   1:   0] slv_grp5_p0_cmd_beat          ;
  wire    [   2:   0] slv_grp5_p0_cmd_usr           ;
  wire                slv_grp5_p0_rsp_ready         ;
  wire                slv_grp5_p0_rsp_valid         ;
  wire                slv_grp5_p0_rsp_err           ;
  wire                slv_grp5_p0_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp5_p0_rsp_rdata         ;
  wire    [   2:   0] slv_grp5_p0_rsp_usr           ;
      wire                slv_grp5_p0_w2n_cmd_valid     ;
  wire                slv_grp5_p0_w2n_cmd_ready     ;
  wire                slv_grp5_p0_w2n_cmd_sel       ;
  wire                slv_grp5_p0_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp5_p0_w2n_cmd_addr      ;
  wire    [  63:   0] slv_grp5_p0_w2n_cmd_wdata     ;
  wire    [   7:   0] slv_grp5_p0_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp5_p0_w2n_cmd_size      ;
  wire                slv_grp5_p0_w2n_cmd_lock      ;
  wire                slv_grp5_p0_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp5_p0_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp5_p0_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp5_p0_w2n_cmd_modes     ;
  wire                slv_grp5_p0_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp5_p0_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp5_p0_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp5_p0_w2n_cmd_usr       ;
  wire                slv_grp5_p0_w2n_rsp_ready     ;
  wire                slv_grp5_p0_w2n_rsp_valid     ;
  wire                slv_grp5_p0_w2n_rsp_err       ;
  wire                slv_grp5_p0_w2n_rsp_excl_ok   ;
  wire    [  63:   0] slv_grp5_p0_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp5_p0_w2n_rsp_usr       ;
      wire                slv_grp5_p0_ro_cmd_valid      ;
  wire                slv_grp5_p0_ro_cmd_ready      ;
  wire                slv_grp5_p0_ro_cmd_sel        ;
  wire                slv_grp5_p0_ro_cmd_read       ;
  wire    [  31:   0] slv_grp5_p0_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp5_p0_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp5_p0_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp5_p0_ro_cmd_size       ;
  wire                slv_grp5_p0_ro_cmd_lock       ;
  wire                slv_grp5_p0_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp5_p0_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp5_p0_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp5_p0_ro_cmd_modes      ;
  wire                slv_grp5_p0_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp5_p0_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp5_p0_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp5_p0_ro_cmd_usr        ;
  wire                slv_grp5_p0_ro_rsp_ready      ;
  wire                slv_grp5_p0_ro_rsp_valid      ;
  wire                slv_grp5_p0_ro_rsp_err        ;
  wire                slv_grp5_p0_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp5_p0_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp5_p0_ro_rsp_usr        ;
      wire                slv_grp5_p0_w2n_ro_cmd_valid  ;
  wire                slv_grp5_p0_w2n_ro_cmd_ready  ;
  wire                slv_grp5_p0_w2n_ro_cmd_sel    ;
  wire                slv_grp5_p0_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp5_p0_w2n_ro_cmd_addr   ;
  wire    [  63:   0] slv_grp5_p0_w2n_ro_cmd_wdata  ;
  wire    [   7:   0] slv_grp5_p0_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp5_p0_w2n_ro_cmd_size   ;
  wire                slv_grp5_p0_w2n_ro_cmd_lock   ;
  wire                slv_grp5_p0_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp5_p0_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp5_p0_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp5_p0_w2n_ro_cmd_modes  ;
  wire                slv_grp5_p0_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp5_p0_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp5_p0_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp5_p0_w2n_ro_cmd_usr    ;
  wire                slv_grp5_p0_w2n_ro_rsp_ready  ;
  wire                slv_grp5_p0_w2n_ro_rsp_valid  ;
  wire                slv_grp5_p0_w2n_ro_rsp_err    ;
  wire                slv_grp5_p0_w2n_ro_rsp_excl_ok ;
  wire    [  63:   0] slv_grp5_p0_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp5_p0_w2n_ro_rsp_usr    ;
      wire                slv_grp5_p0_wo_cmd_valid      ;
  wire                slv_grp5_p0_wo_cmd_ready      ;
  wire                slv_grp5_p0_wo_cmd_sel        ;
  wire                slv_grp5_p0_wo_cmd_read       ;
  wire    [  31:   0] slv_grp5_p0_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp5_p0_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp5_p0_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp5_p0_wo_cmd_size       ;
  wire                slv_grp5_p0_wo_cmd_lock       ;
  wire                slv_grp5_p0_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp5_p0_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp5_p0_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp5_p0_wo_cmd_modes      ;
  wire                slv_grp5_p0_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp5_p0_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp5_p0_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp5_p0_wo_cmd_usr        ;
  wire                slv_grp5_p0_wo_rsp_ready      ;
  wire                slv_grp5_p0_wo_rsp_valid      ;
  wire                slv_grp5_p0_wo_rsp_err        ;
  wire                slv_grp5_p0_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp5_p0_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp5_p0_wo_rsp_usr        ;
      wire                slv_grp5_p0_w2n_wo_cmd_valid  ;
  wire                slv_grp5_p0_w2n_wo_cmd_ready  ;
  wire                slv_grp5_p0_w2n_wo_cmd_sel    ;
  wire                slv_grp5_p0_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp5_p0_w2n_wo_cmd_addr   ;
  wire    [  63:   0] slv_grp5_p0_w2n_wo_cmd_wdata  ;
  wire    [   7:   0] slv_grp5_p0_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp5_p0_w2n_wo_cmd_size   ;
  wire                slv_grp5_p0_w2n_wo_cmd_lock   ;
  wire                slv_grp5_p0_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp5_p0_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp5_p0_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp5_p0_w2n_wo_cmd_modes  ;
  wire                slv_grp5_p0_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp5_p0_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp5_p0_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp5_p0_w2n_wo_cmd_usr    ;
  wire                slv_grp5_p0_w2n_wo_rsp_ready  ;
  wire                slv_grp5_p0_w2n_wo_rsp_valid  ;
  wire                slv_grp5_p0_w2n_wo_rsp_err    ;
  wire                slv_grp5_p0_w2n_wo_rsp_excl_ok ;
  wire    [  63:   0] slv_grp5_p0_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp5_p0_w2n_wo_rsp_usr    ;
                wire                      slv_grp5_p0_w2n_wo_rsp_last;
   e603_subsys_sgrp5_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (32'h80000000),
      .O0_BASE_REGION_LSB(31),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (128 ),
      .SPLT_FIFO_OUTS_CNT_W(8),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp5_ro_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_5_ro_icb_cmd_valid               ),
  .i_icb_cmd_ready                (slv_grp_5_ro_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (slv_grp_5_ro_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (slv_grp_5_ro_icb_cmd_read                ),
  .i_icb_cmd_addr                 (slv_grp_5_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_5_ro_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_5_ro_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_5_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_5_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (slv_grp_5_ro_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (slv_grp_5_ro_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_5_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_5_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_5_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (slv_grp_5_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_5_ro_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_5_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_5_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (slv_grp_5_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (slv_grp_5_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (slv_grp_5_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (slv_grp_5_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_5_ro_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (slv_grp5_p0_ro_cmd_valid                 ),
  .o0_icb_cmd_ready               (slv_grp5_p0_ro_cmd_ready                 ),
  .o0_icb_cmd_sel                 (slv_grp5_p0_ro_cmd_sel                   ),
  .o0_icb_cmd_read                (slv_grp5_p0_ro_cmd_read                  ),
  .o0_icb_cmd_addr                (slv_grp5_p0_ro_cmd_addr       [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp5_p0_ro_cmd_wdata      [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp5_p0_ro_cmd_wmask      [   7:   0]),
  .o0_icb_cmd_size                (slv_grp5_p0_ro_cmd_size       [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp5_p0_ro_cmd_lock                  ),
  .o0_icb_cmd_excl                (slv_grp5_p0_ro_cmd_excl                  ),
  .o0_icb_cmd_xlen                (slv_grp5_p0_ro_cmd_xlen       [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp5_p0_ro_cmd_xburst     [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp5_p0_ro_cmd_modes      [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp5_p0_ro_cmd_dmode                 ),
  .o0_icb_cmd_attri               (slv_grp5_p0_ro_cmd_attri      [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp5_p0_ro_cmd_beat       [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp5_p0_ro_cmd_usr        [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp5_p0_ro_rsp_ready                 ),
  .o0_icb_rsp_valid               (slv_grp5_p0_ro_rsp_valid                 ),
  .o0_icb_rsp_err                 (slv_grp5_p0_ro_rsp_err                   ),
  .o0_icb_rsp_excl_ok             (slv_grp5_p0_ro_rsp_excl_ok               ),
  .o0_icb_rsp_rdata               (slv_grp5_p0_ro_rsp_rdata      [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp5_p0_ro_rsp_usr        [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_sgrp5_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (0),
      .ICB_FIFO_CMD_DP        (2),
      .ICB_FIFO_RSP_DP        (2),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (32'h80000000),
      .O0_BASE_REGION_LSB(31),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (128 ),
      .SPLT_FIFO_OUTS_CNT_W(8),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp5_wo_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_5_wo_icb_cmd_valid               ),
  .i_icb_cmd_ready                (slv_grp_5_wo_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (slv_grp_5_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (slv_grp_5_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (slv_grp_5_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_5_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_5_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_5_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_5_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (slv_grp_5_wo_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (slv_grp_5_wo_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_5_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_5_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_5_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (slv_grp_5_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_5_wo_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_5_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_5_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (slv_grp_5_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (slv_grp_5_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (slv_grp_5_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (slv_grp_5_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_5_wo_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (slv_grp5_p0_wo_cmd_valid                 ),
  .o0_icb_cmd_ready               (slv_grp5_p0_wo_cmd_ready                 ),
  .o0_icb_cmd_sel                 (slv_grp5_p0_wo_cmd_sel                   ),
  .o0_icb_cmd_read                (slv_grp5_p0_wo_cmd_read                  ),
  .o0_icb_cmd_addr                (slv_grp5_p0_wo_cmd_addr       [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp5_p0_wo_cmd_wdata      [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp5_p0_wo_cmd_wmask      [   7:   0]),
  .o0_icb_cmd_size                (slv_grp5_p0_wo_cmd_size       [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp5_p0_wo_cmd_lock                  ),
  .o0_icb_cmd_excl                (slv_grp5_p0_wo_cmd_excl                  ),
  .o0_icb_cmd_xlen                (slv_grp5_p0_wo_cmd_xlen       [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp5_p0_wo_cmd_xburst     [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp5_p0_wo_cmd_modes      [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp5_p0_wo_cmd_dmode                 ),
  .o0_icb_cmd_attri               (slv_grp5_p0_wo_cmd_attri      [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp5_p0_wo_cmd_beat       [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp5_p0_wo_cmd_usr        [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp5_p0_wo_rsp_ready                 ),
  .o0_icb_rsp_valid               (slv_grp5_p0_wo_rsp_valid                 ),
  .o0_icb_rsp_err                 (slv_grp5_p0_wo_rsp_err                   ),
  .o0_icb_rsp_excl_ok             (slv_grp5_p0_wo_rsp_excl_ok               ),
  .o0_icb_rsp_rdata               (slv_grp5_p0_wo_rsp_rdata      [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp5_p0_wo_rsp_usr        [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (128),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_o0_axi_ro_icb_wconv(
      .i_icb_cmd_read(1'b1),
      .i_icb_cmd_wdata(64'b0),
      .i_icb_cmd_wmask(8'b0),
        .i_icb_cmd_valid                (slv_grp5_p0_ro_cmd_valid                 ),
  .i_icb_cmd_ready                (slv_grp5_p0_ro_cmd_ready                 ),
  .i_icb_cmd_sel                  (slv_grp5_p0_ro_cmd_sel                   ),
  .i_icb_cmd_addr                 (slv_grp5_p0_ro_cmd_addr       [  31:   0]),
  .i_icb_cmd_size                 (slv_grp5_p0_ro_cmd_size       [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp5_p0_ro_cmd_lock                  ),
  .i_icb_cmd_excl                 (slv_grp5_p0_ro_cmd_excl                  ),
  .i_icb_cmd_xlen                 (slv_grp5_p0_ro_cmd_xlen       [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp5_p0_ro_cmd_xburst     [   1:   0]),
  .i_icb_cmd_modes                (slv_grp5_p0_ro_cmd_modes      [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp5_p0_ro_cmd_dmode                 ),
  .i_icb_cmd_attri                (slv_grp5_p0_ro_cmd_attri      [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp5_p0_ro_cmd_beat       [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp5_p0_ro_cmd_usr        [   2:   0]),
  .i_icb_rsp_ready                (slv_grp5_p0_ro_rsp_ready                 ),
  .i_icb_rsp_valid                (slv_grp5_p0_ro_rsp_valid                 ),
  .i_icb_rsp_err                  (slv_grp5_p0_ro_rsp_err                   ),
  .i_icb_rsp_excl_ok              (slv_grp5_p0_ro_rsp_excl_ok               ),
  .i_icb_rsp_rdata                (slv_grp5_p0_ro_rsp_rdata      [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp5_p0_ro_rsp_usr        [   2:   0]),
        .o_icb_cmd_valid                (slv_grp5_p0_w2n_ro_cmd_valid             ),
  .o_icb_cmd_ready                (slv_grp5_p0_w2n_ro_cmd_ready             ),
  .o_icb_cmd_sel                  (slv_grp5_p0_w2n_ro_cmd_sel               ),
  .o_icb_cmd_read                 (slv_grp5_p0_w2n_ro_cmd_read              ),
  .o_icb_cmd_addr                 (slv_grp5_p0_w2n_ro_cmd_addr   [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp5_p0_w2n_ro_cmd_wdata  [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp5_p0_w2n_ro_cmd_wmask  [   7:   0]),
  .o_icb_cmd_size                 (slv_grp5_p0_w2n_ro_cmd_size   [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp5_p0_w2n_ro_cmd_lock              ),
  .o_icb_cmd_excl                 (slv_grp5_p0_w2n_ro_cmd_excl              ),
  .o_icb_cmd_xlen                 (slv_grp5_p0_w2n_ro_cmd_xlen   [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp5_p0_w2n_ro_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (slv_grp5_p0_w2n_ro_cmd_modes  [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp5_p0_w2n_ro_cmd_dmode             ),
  .o_icb_cmd_attri                (slv_grp5_p0_w2n_ro_cmd_attri  [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp5_p0_w2n_ro_cmd_beat   [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp5_p0_w2n_ro_cmd_usr    [   2:   0]),
  .o_icb_rsp_ready                (slv_grp5_p0_w2n_ro_rsp_ready             ),
  .o_icb_rsp_valid                (slv_grp5_p0_w2n_ro_rsp_valid             ),
  .o_icb_rsp_err                  (slv_grp5_p0_w2n_ro_rsp_err               ),
  .o_icb_rsp_excl_ok              (slv_grp5_p0_w2n_ro_rsp_excl_ok            ),
  .o_icb_rsp_rdata                (slv_grp5_p0_w2n_ro_rsp_rdata  [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp5_p0_w2n_ro_rsp_usr    [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (128),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_o0_axi_wo_icb_wconv(
        .i_icb_cmd_valid                (slv_grp5_p0_wo_cmd_valid                 ),
  .i_icb_cmd_ready                (slv_grp5_p0_wo_cmd_ready                 ),
  .i_icb_cmd_sel                  (slv_grp5_p0_wo_cmd_sel                   ),
  .i_icb_cmd_read                 (slv_grp5_p0_wo_cmd_read                  ),
  .i_icb_cmd_addr                 (slv_grp5_p0_wo_cmd_addr       [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp5_p0_wo_cmd_wdata      [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp5_p0_wo_cmd_wmask      [   7:   0]),
  .i_icb_cmd_size                 (slv_grp5_p0_wo_cmd_size       [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp5_p0_wo_cmd_lock                  ),
  .i_icb_cmd_excl                 (slv_grp5_p0_wo_cmd_excl                  ),
  .i_icb_cmd_xlen                 (slv_grp5_p0_wo_cmd_xlen       [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp5_p0_wo_cmd_xburst     [   1:   0]),
  .i_icb_cmd_modes                (slv_grp5_p0_wo_cmd_modes      [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp5_p0_wo_cmd_dmode                 ),
  .i_icb_cmd_attri                (slv_grp5_p0_wo_cmd_attri      [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp5_p0_wo_cmd_beat       [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp5_p0_wo_cmd_usr        [   2:   0]),
  .i_icb_rsp_ready                (slv_grp5_p0_wo_rsp_ready                 ),
  .i_icb_rsp_valid                (slv_grp5_p0_wo_rsp_valid                 ),
  .i_icb_rsp_err                  (slv_grp5_p0_wo_rsp_err                   ),
  .i_icb_rsp_excl_ok              (slv_grp5_p0_wo_rsp_excl_ok               ),
  .i_icb_rsp_rdata                (slv_grp5_p0_wo_rsp_rdata      [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp5_p0_wo_rsp_usr        [   2:   0]),
      .o_icb_rsp_rdata(64'b0),
        .o_icb_cmd_valid                (slv_grp5_p0_w2n_wo_cmd_valid             ),
  .o_icb_cmd_ready                (slv_grp5_p0_w2n_wo_cmd_ready             ),
  .o_icb_cmd_sel                  (slv_grp5_p0_w2n_wo_cmd_sel               ),
  .o_icb_cmd_read                 (slv_grp5_p0_w2n_wo_cmd_read              ),
  .o_icb_cmd_addr                 (slv_grp5_p0_w2n_wo_cmd_addr   [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp5_p0_w2n_wo_cmd_wdata  [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp5_p0_w2n_wo_cmd_wmask  [   7:   0]),
  .o_icb_cmd_size                 (slv_grp5_p0_w2n_wo_cmd_size   [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp5_p0_w2n_wo_cmd_lock              ),
  .o_icb_cmd_excl                 (slv_grp5_p0_w2n_wo_cmd_excl              ),
  .o_icb_cmd_xlen                 (slv_grp5_p0_w2n_wo_cmd_xlen   [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp5_p0_w2n_wo_cmd_xburst [   1:   0]),
  .o_icb_cmd_modes                (slv_grp5_p0_w2n_wo_cmd_modes  [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp5_p0_w2n_wo_cmd_dmode             ),
  .o_icb_cmd_attri                (slv_grp5_p0_w2n_wo_cmd_attri  [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp5_p0_w2n_wo_cmd_beat   [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp5_p0_w2n_wo_cmd_usr    [   2:   0]),
  .o_icb_rsp_ready                (slv_grp5_p0_w2n_wo_rsp_ready             ),
  .o_icb_rsp_valid                (slv_grp5_p0_w2n_wo_rsp_valid             ),
  .o_icb_rsp_err                  (slv_grp5_p0_w2n_wo_rsp_err               ),
  .o_icb_rsp_excl_ok              (slv_grp5_p0_w2n_wo_rsp_excl_ok            ),
  .o_icb_rsp_usr                  (slv_grp5_p0_w2n_wo_rsp_usr    [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      wire o0_axi_ro_bus_pend_active;
      wire o0_axi_ro_bus_icb_active;
      wire o0_axi_wo_bus_pend_active;
      wire o0_axi_wo_bus_icb_active;
      wire o0_axi_bus_pend_active = 1'b0 
                                   | o0_axi_ro_bus_pend_active 
                                   | o0_axi_wo_bus_pend_active
                                   ;
      wire o0_axi_bus_icb_active = 1'b0 
                                   | o0_axi_ro_bus_icb_active 
                                   | o0_axi_wo_bus_icb_active
                                   ;
      assign o0_axi_arid = 3'b0;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(8+1)
      )u_o0_axi__ro_icb_active (
         .icb_active(o0_axi_ro_bus_icb_active),
            .icb_cmd_valid(slv_grp5_p0_w2n_ro_cmd_valid),
            .icb_cmd_ready(slv_grp5_p0_w2n_ro_cmd_ready),
            .icb_rsp_valid(slv_grp5_p0_w2n_ro_rsp_valid),
            .icb_rsp_ready(slv_grp5_p0_w2n_ro_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] o0_axi_araddr_full;
      assign o0_axi_araddr = o0_axi_araddr_full[32-1:0];
  e603_subsys_gnrl_ficb2axi_read_async # (
    .SYNC_DP       (2),
    .ASYNC_FIFO    (1),
    .ASYNC_FIFO_DP (8),
    .ASYNC_FIFO_DP_PTR_W (3),
    .AW    (32),
    .DW    (64),
    .OUTS_CNT_W (8 ),
    .CMD_UW (3),
    .RSP_UW (3)
    ) u_o0_axi_icb2axi_read(
    .icb2axi_read_pend_active(o0_axi_ro_bus_pend_active),
      .icb_cmd_valid                  (slv_grp5_p0_w2n_ro_cmd_valid             ),
  .icb_cmd_ready                  (slv_grp5_p0_w2n_ro_cmd_ready             ),
  .icb_cmd_sel                    (slv_grp5_p0_w2n_ro_cmd_sel               ),
  .icb_cmd_read                   (slv_grp5_p0_w2n_ro_cmd_read              ),
  .icb_cmd_wdata                  (slv_grp5_p0_w2n_ro_cmd_wdata  [  63:   0]),
  .icb_cmd_wmask                  (slv_grp5_p0_w2n_ro_cmd_wmask  [   7:   0]),
  .icb_cmd_size                   (slv_grp5_p0_w2n_ro_cmd_size   [   2:   0]),
  .icb_cmd_lock                   (slv_grp5_p0_w2n_ro_cmd_lock              ),
  .icb_cmd_excl                   (slv_grp5_p0_w2n_ro_cmd_excl              ),
  .icb_cmd_xlen                   (slv_grp5_p0_w2n_ro_cmd_xlen   [   7:   0]),
  .icb_cmd_xburst                 (slv_grp5_p0_w2n_ro_cmd_xburst [   1:   0]),
  .icb_cmd_modes                  (slv_grp5_p0_w2n_ro_cmd_modes  [   1:   0]),
  .icb_cmd_dmode                  (slv_grp5_p0_w2n_ro_cmd_dmode             ),
  .icb_cmd_attri                  (slv_grp5_p0_w2n_ro_cmd_attri  [   2:   0]),
  .icb_cmd_beat                   (slv_grp5_p0_w2n_ro_cmd_beat   [   1:   0]),
  .icb_rsp_ready                  (slv_grp5_p0_w2n_ro_rsp_ready             ),
  .icb_rsp_valid                  (slv_grp5_p0_w2n_ro_rsp_valid             ),
  .icb_rsp_err                    (slv_grp5_p0_w2n_ro_rsp_err               ),
  .icb_rsp_excl_ok                (slv_grp5_p0_w2n_ro_rsp_excl_ok            ),
  .icb_rsp_rdata                  (slv_grp5_p0_w2n_ro_rsp_rdata  [  63:   0]),
             .icb_cmd_usr(slv_grp5_p0_w2n_ro_cmd_usr[3-1:0]),
             .icb_rsp_usr(slv_grp5_p0_w2n_ro_rsp_usr[3-1:0]),
      .icb_cmd_addr(slv_grp5_p0_w2n_ro_cmd_addr),
      .axi_araddr(o0_axi_araddr_full),
      .axi_arvalid                    (o0_axi_arvalid                           ),
  .axi_arready                    (o0_axi_arready                           ),
  .axi_arlen                      (o0_axi_arlen                  [   7:   0]),
  .axi_arsize                     (o0_axi_arsize                 [   2:   0]),
  .axi_arburst                    (o0_axi_arburst                [   1:   0]),
  .axi_arlock                     (o0_axi_arlock                            ),
  .axi_arcache                    (o0_axi_arcache                [   3:   0]),
  .axi_arprot                     (o0_axi_arprot                 [   2:   0]),
  .axi_rready                     (o0_axi_rready                            ),
  .axi_rvalid                     (o0_axi_rvalid                            ),
  .axi_rdata                      (o0_axi_rdata                  [  63:   0]),
  .axi_rresp                      (o0_axi_rresp                  [   1:   0]),
  .axi_rlast                      (o0_axi_rlast                             ),
      .axi_aruser(),
      .axi_ruser(3'b0),
    .icb2axi_read_async_icb_active(),
    .icb2axi_read_async_axi_active(),
    .async_axi_clk  (o0_axi_clk  ),
    .async_axi_rst_n(o0_axi_rst_n_sync_4port),
    .icb_clk        (clk),
    .icb_rst_n      (o0_axi_rst_n_sync_4fab)
  );
       assign o0_axi_awid = 3'b0;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(8+1)
      )u_o0_axi__wo_icb_active (
         .icb_active(o0_axi_wo_bus_icb_active),
            .icb_cmd_valid(slv_grp5_p0_w2n_wo_cmd_valid),
            .icb_cmd_ready(slv_grp5_p0_w2n_wo_cmd_ready),
            .icb_rsp_valid(slv_grp5_p0_w2n_wo_rsp_valid),
            .icb_rsp_ready(slv_grp5_p0_w2n_wo_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] o0_axi_awaddr_full;
      assign o0_axi_awaddr = o0_axi_awaddr_full[32-1:0];
  e603_subsys_gnrl_ficb2axi_write_async # (
    .SYNC_DP       (2),
    .ASYNC_FIFO    (1),
    .ASYNC_FIFO_DP (8),
    .ASYNC_FIFO_DP_PTR_W (3),
    .AW    (32),
    .DW    (64),
    .OUTS_FIFO_DP (128 ),
    .OUTS_CNT_W (8 ),
    .CMD_UW (3),
    .RSP_UW (3)
    ) u_o0_axi_icb2axi_write(
    .icb2axi_write_pend_active(o0_axi_wo_bus_pend_active),
      .icb_cmd_valid                  (slv_grp5_p0_w2n_wo_cmd_valid             ),
  .icb_cmd_ready                  (slv_grp5_p0_w2n_wo_cmd_ready             ),
  .icb_cmd_sel                    (slv_grp5_p0_w2n_wo_cmd_sel               ),
  .icb_cmd_read                   (slv_grp5_p0_w2n_wo_cmd_read              ),
  .icb_cmd_wdata                  (slv_grp5_p0_w2n_wo_cmd_wdata  [  63:   0]),
  .icb_cmd_wmask                  (slv_grp5_p0_w2n_wo_cmd_wmask  [   7:   0]),
  .icb_cmd_size                   (slv_grp5_p0_w2n_wo_cmd_size   [   2:   0]),
  .icb_cmd_lock                   (slv_grp5_p0_w2n_wo_cmd_lock              ),
  .icb_cmd_excl                   (slv_grp5_p0_w2n_wo_cmd_excl              ),
  .icb_cmd_xlen                   (slv_grp5_p0_w2n_wo_cmd_xlen   [   7:   0]),
  .icb_cmd_xburst                 (slv_grp5_p0_w2n_wo_cmd_xburst [   1:   0]),
  .icb_cmd_modes                  (slv_grp5_p0_w2n_wo_cmd_modes  [   1:   0]),
  .icb_cmd_dmode                  (slv_grp5_p0_w2n_wo_cmd_dmode             ),
  .icb_cmd_attri                  (slv_grp5_p0_w2n_wo_cmd_attri  [   2:   0]),
  .icb_cmd_beat                   (slv_grp5_p0_w2n_wo_cmd_beat   [   1:   0]),
  .icb_rsp_ready                  (slv_grp5_p0_w2n_wo_rsp_ready             ),
  .icb_rsp_valid                  (slv_grp5_p0_w2n_wo_rsp_valid             ),
  .icb_rsp_err                    (slv_grp5_p0_w2n_wo_rsp_err               ),
  .icb_rsp_excl_ok                (slv_grp5_p0_w2n_wo_rsp_excl_ok            ),
  .icb_rsp_rdata                  (slv_grp5_p0_w2n_wo_rsp_rdata  [  63:   0]),
             .icb_cmd_usr(slv_grp5_p0_w2n_wo_cmd_usr[3-1:0]),
             .icb_rsp_usr(slv_grp5_p0_w2n_wo_rsp_usr[3-1:0]),
      .icb_cmd_addr(slv_grp5_p0_w2n_wo_cmd_addr),
      .axi_awaddr(o0_axi_awaddr_full),
      .axi_awvalid                    (o0_axi_awvalid                           ),
  .axi_awready                    (o0_axi_awready                           ),
  .axi_awlen                      (o0_axi_awlen                  [   7:   0]),
  .axi_awsize                     (o0_axi_awsize                 [   2:   0]),
  .axi_awburst                    (o0_axi_awburst                [   1:   0]),
  .axi_awlock                     (o0_axi_awlock                            ),
  .axi_awcache                    (o0_axi_awcache                [   3:   0]),
  .axi_awprot                     (o0_axi_awprot                 [   2:   0]),
  .axi_bready                     (o0_axi_bready                            ),
  .axi_bvalid                     (o0_axi_bvalid                            ),
  .axi_bresp                      (o0_axi_bresp                  [   1:   0]),
  .axi_wready                     (o0_axi_wready                            ),
  .axi_wvalid                     (o0_axi_wvalid                            ),
  .axi_wdata                      (o0_axi_wdata                  [  63:   0]),
  .axi_wstrb                      (o0_axi_wstrb                  [   7:   0]),
  .axi_wlast                      (o0_axi_wlast                             ),
      .axi_awuser(),
      .axi_buser(3'b0),
    .icb2axi_write_async_icb_active(),
    .icb2axi_write_async_axi_active(),
    .async_axi_clk  (o0_axi_clk  ),
    .async_axi_rst_n(o0_axi_rst_n_sync_4port),
    .icb_clk        (clk),
    .icb_rst_n      (o0_axi_rst_n_sync_4fab)
  );
      wire                slv_grp_6_icb_cmd_valid       ;
  wire                slv_grp_6_icb_cmd_ready       ;
  wire                slv_grp_6_icb_cmd_sel         ;
  wire                slv_grp_6_icb_cmd_read        ;
  wire    [  31:   0] slv_grp_6_icb_cmd_addr        ;
  wire    [  63:   0] slv_grp_6_icb_cmd_wdata       ;
  wire    [   7:   0] slv_grp_6_icb_cmd_wmask       ;
  wire    [   2:   0] slv_grp_6_icb_cmd_size        ;
  wire                slv_grp_6_icb_cmd_lock        ;
  wire                slv_grp_6_icb_cmd_excl        ;
  wire    [   7:   0] slv_grp_6_icb_cmd_xlen        ;
  wire    [   1:   0] slv_grp_6_icb_cmd_xburst      ;
  wire    [   1:   0] slv_grp_6_icb_cmd_modes       ;
  wire                slv_grp_6_icb_cmd_dmode       ;
  wire    [   2:   0] slv_grp_6_icb_cmd_attri       ;
  wire    [   1:   0] slv_grp_6_icb_cmd_beat        ;
  wire    [   2:   0] slv_grp_6_icb_cmd_usr         ;
  wire                slv_grp_6_icb_rsp_ready       ;
  wire                slv_grp_6_icb_rsp_valid       ;
  wire                slv_grp_6_icb_rsp_err         ;
  wire                slv_grp_6_icb_rsp_excl_ok     ;
  wire    [  63:   0] slv_grp_6_icb_rsp_rdata       ;
  wire    [   2:   0] slv_grp_6_icb_rsp_usr         ;
      wire                slv_grp_6_ro_icb_cmd_valid    ;
  wire                slv_grp_6_ro_icb_cmd_ready    ;
  wire                slv_grp_6_ro_icb_cmd_sel      ;
  wire                slv_grp_6_ro_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_6_ro_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_6_ro_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_6_ro_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_6_ro_icb_cmd_size     ;
  wire                slv_grp_6_ro_icb_cmd_lock     ;
  wire                slv_grp_6_ro_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_6_ro_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_6_ro_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_6_ro_icb_cmd_modes    ;
  wire                slv_grp_6_ro_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_6_ro_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_6_ro_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_6_ro_icb_cmd_usr      ;
  wire                slv_grp_6_ro_icb_rsp_ready    ;
  wire                slv_grp_6_ro_icb_rsp_valid    ;
  wire                slv_grp_6_ro_icb_rsp_err      ;
  wire                slv_grp_6_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_6_ro_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_6_ro_icb_rsp_usr      ;
      wire                slv_grp_6_wo_icb_cmd_valid    ;
  wire                slv_grp_6_wo_icb_cmd_ready    ;
  wire                slv_grp_6_wo_icb_cmd_sel      ;
  wire                slv_grp_6_wo_icb_cmd_read     ;
  wire    [  31:   0] slv_grp_6_wo_icb_cmd_addr     ;
  wire    [  63:   0] slv_grp_6_wo_icb_cmd_wdata    ;
  wire    [   7:   0] slv_grp_6_wo_icb_cmd_wmask    ;
  wire    [   2:   0] slv_grp_6_wo_icb_cmd_size     ;
  wire                slv_grp_6_wo_icb_cmd_lock     ;
  wire                slv_grp_6_wo_icb_cmd_excl     ;
  wire    [   7:   0] slv_grp_6_wo_icb_cmd_xlen     ;
  wire    [   1:   0] slv_grp_6_wo_icb_cmd_xburst   ;
  wire    [   1:   0] slv_grp_6_wo_icb_cmd_modes    ;
  wire                slv_grp_6_wo_icb_cmd_dmode    ;
  wire    [   2:   0] slv_grp_6_wo_icb_cmd_attri    ;
  wire    [   1:   0] slv_grp_6_wo_icb_cmd_beat     ;
  wire    [   2:   0] slv_grp_6_wo_icb_cmd_usr      ;
  wire                slv_grp_6_wo_icb_rsp_ready    ;
  wire                slv_grp_6_wo_icb_rsp_valid    ;
  wire                slv_grp_6_wo_icb_rsp_err      ;
  wire                slv_grp_6_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] slv_grp_6_wo_icb_rsp_rdata    ;
  wire    [   2:   0] slv_grp_6_wo_icb_rsp_usr      ;
      wire                slv_grp6_p0_cmd_valid         ;
  wire                slv_grp6_p0_cmd_ready         ;
  wire                slv_grp6_p0_cmd_sel           ;
  wire                slv_grp6_p0_cmd_read          ;
  wire    [  31:   0] slv_grp6_p0_cmd_addr          ;
  wire    [  63:   0] slv_grp6_p0_cmd_wdata         ;
  wire    [   7:   0] slv_grp6_p0_cmd_wmask         ;
  wire    [   2:   0] slv_grp6_p0_cmd_size          ;
  wire                slv_grp6_p0_cmd_lock          ;
  wire                slv_grp6_p0_cmd_excl          ;
  wire    [   7:   0] slv_grp6_p0_cmd_xlen          ;
  wire    [   1:   0] slv_grp6_p0_cmd_xburst        ;
  wire    [   1:   0] slv_grp6_p0_cmd_modes         ;
  wire                slv_grp6_p0_cmd_dmode         ;
  wire    [   2:   0] slv_grp6_p0_cmd_attri         ;
  wire    [   1:   0] slv_grp6_p0_cmd_beat          ;
  wire    [   2:   0] slv_grp6_p0_cmd_usr           ;
  wire                slv_grp6_p0_rsp_ready         ;
  wire                slv_grp6_p0_rsp_valid         ;
  wire                slv_grp6_p0_rsp_err           ;
  wire                slv_grp6_p0_rsp_excl_ok       ;
  wire    [  63:   0] slv_grp6_p0_rsp_rdata         ;
  wire    [   2:   0] slv_grp6_p0_rsp_usr           ;
      wire                slv_grp6_p0_w2n_cmd_valid     ;
  wire                slv_grp6_p0_w2n_cmd_ready     ;
  wire                slv_grp6_p0_w2n_cmd_sel       ;
  wire                slv_grp6_p0_w2n_cmd_read      ;
  wire    [  31:   0] slv_grp6_p0_w2n_cmd_addr      ;
  wire    [  63:   0] slv_grp6_p0_w2n_cmd_wdata     ;
  wire    [   7:   0] slv_grp6_p0_w2n_cmd_wmask     ;
  wire    [   2:   0] slv_grp6_p0_w2n_cmd_size      ;
  wire                slv_grp6_p0_w2n_cmd_lock      ;
  wire                slv_grp6_p0_w2n_cmd_excl      ;
  wire    [   7:   0] slv_grp6_p0_w2n_cmd_xlen      ;
  wire    [   1:   0] slv_grp6_p0_w2n_cmd_xburst    ;
  wire    [   1:   0] slv_grp6_p0_w2n_cmd_modes     ;
  wire                slv_grp6_p0_w2n_cmd_dmode     ;
  wire    [   2:   0] slv_grp6_p0_w2n_cmd_attri     ;
  wire    [   1:   0] slv_grp6_p0_w2n_cmd_beat      ;
  wire    [   2:   0] slv_grp6_p0_w2n_cmd_usr       ;
  wire                slv_grp6_p0_w2n_rsp_ready     ;
  wire                slv_grp6_p0_w2n_rsp_valid     ;
  wire                slv_grp6_p0_w2n_rsp_err       ;
  wire                slv_grp6_p0_w2n_rsp_excl_ok   ;
  wire    [  63:   0] slv_grp6_p0_w2n_rsp_rdata     ;
  wire    [   2:   0] slv_grp6_p0_w2n_rsp_usr       ;
      wire                slv_grp6_p0_ro_cmd_valid      ;
  wire                slv_grp6_p0_ro_cmd_ready      ;
  wire                slv_grp6_p0_ro_cmd_sel        ;
  wire                slv_grp6_p0_ro_cmd_read       ;
  wire    [  31:   0] slv_grp6_p0_ro_cmd_addr       ;
  wire    [  63:   0] slv_grp6_p0_ro_cmd_wdata      ;
  wire    [   7:   0] slv_grp6_p0_ro_cmd_wmask      ;
  wire    [   2:   0] slv_grp6_p0_ro_cmd_size       ;
  wire                slv_grp6_p0_ro_cmd_lock       ;
  wire                slv_grp6_p0_ro_cmd_excl       ;
  wire    [   7:   0] slv_grp6_p0_ro_cmd_xlen       ;
  wire    [   1:   0] slv_grp6_p0_ro_cmd_xburst     ;
  wire    [   1:   0] slv_grp6_p0_ro_cmd_modes      ;
  wire                slv_grp6_p0_ro_cmd_dmode      ;
  wire    [   2:   0] slv_grp6_p0_ro_cmd_attri      ;
  wire    [   1:   0] slv_grp6_p0_ro_cmd_beat       ;
  wire    [   2:   0] slv_grp6_p0_ro_cmd_usr        ;
  wire                slv_grp6_p0_ro_rsp_ready      ;
  wire                slv_grp6_p0_ro_rsp_valid      ;
  wire                slv_grp6_p0_ro_rsp_err        ;
  wire                slv_grp6_p0_ro_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp6_p0_ro_rsp_rdata      ;
  wire    [   2:   0] slv_grp6_p0_ro_rsp_usr        ;
      wire                slv_grp6_p0_w2n_ro_cmd_valid  ;
  wire                slv_grp6_p0_w2n_ro_cmd_ready  ;
  wire                slv_grp6_p0_w2n_ro_cmd_sel    ;
  wire                slv_grp6_p0_w2n_ro_cmd_read   ;
  wire    [  31:   0] slv_grp6_p0_w2n_ro_cmd_addr   ;
  wire    [  63:   0] slv_grp6_p0_w2n_ro_cmd_wdata  ;
  wire    [   7:   0] slv_grp6_p0_w2n_ro_cmd_wmask  ;
  wire    [   2:   0] slv_grp6_p0_w2n_ro_cmd_size   ;
  wire                slv_grp6_p0_w2n_ro_cmd_lock   ;
  wire                slv_grp6_p0_w2n_ro_cmd_excl   ;
  wire    [   7:   0] slv_grp6_p0_w2n_ro_cmd_xlen   ;
  wire    [   1:   0] slv_grp6_p0_w2n_ro_cmd_xburst ;
  wire    [   1:   0] slv_grp6_p0_w2n_ro_cmd_modes  ;
  wire                slv_grp6_p0_w2n_ro_cmd_dmode  ;
  wire    [   2:   0] slv_grp6_p0_w2n_ro_cmd_attri  ;
  wire    [   1:   0] slv_grp6_p0_w2n_ro_cmd_beat   ;
  wire    [   2:   0] slv_grp6_p0_w2n_ro_cmd_usr    ;
  wire                slv_grp6_p0_w2n_ro_rsp_ready  ;
  wire                slv_grp6_p0_w2n_ro_rsp_valid  ;
  wire                slv_grp6_p0_w2n_ro_rsp_err    ;
  wire                slv_grp6_p0_w2n_ro_rsp_excl_ok ;
  wire    [  63:   0] slv_grp6_p0_w2n_ro_rsp_rdata  ;
  wire    [   2:   0] slv_grp6_p0_w2n_ro_rsp_usr    ;
      wire                slv_grp6_p0_wo_cmd_valid      ;
  wire                slv_grp6_p0_wo_cmd_ready      ;
  wire                slv_grp6_p0_wo_cmd_sel        ;
  wire                slv_grp6_p0_wo_cmd_read       ;
  wire    [  31:   0] slv_grp6_p0_wo_cmd_addr       ;
  wire    [  63:   0] slv_grp6_p0_wo_cmd_wdata      ;
  wire    [   7:   0] slv_grp6_p0_wo_cmd_wmask      ;
  wire    [   2:   0] slv_grp6_p0_wo_cmd_size       ;
  wire                slv_grp6_p0_wo_cmd_lock       ;
  wire                slv_grp6_p0_wo_cmd_excl       ;
  wire    [   7:   0] slv_grp6_p0_wo_cmd_xlen       ;
  wire    [   1:   0] slv_grp6_p0_wo_cmd_xburst     ;
  wire    [   1:   0] slv_grp6_p0_wo_cmd_modes      ;
  wire                slv_grp6_p0_wo_cmd_dmode      ;
  wire    [   2:   0] slv_grp6_p0_wo_cmd_attri      ;
  wire    [   1:   0] slv_grp6_p0_wo_cmd_beat       ;
  wire    [   2:   0] slv_grp6_p0_wo_cmd_usr        ;
  wire                slv_grp6_p0_wo_rsp_ready      ;
  wire                slv_grp6_p0_wo_rsp_valid      ;
  wire                slv_grp6_p0_wo_rsp_err        ;
  wire                slv_grp6_p0_wo_rsp_excl_ok    ;
  wire    [  63:   0] slv_grp6_p0_wo_rsp_rdata      ;
  wire    [   2:   0] slv_grp6_p0_wo_rsp_usr        ;
      wire                slv_grp6_p0_w2n_wo_cmd_valid  ;
  wire                slv_grp6_p0_w2n_wo_cmd_ready  ;
  wire                slv_grp6_p0_w2n_wo_cmd_sel    ;
  wire                slv_grp6_p0_w2n_wo_cmd_read   ;
  wire    [  31:   0] slv_grp6_p0_w2n_wo_cmd_addr   ;
  wire    [  63:   0] slv_grp6_p0_w2n_wo_cmd_wdata  ;
  wire    [   7:   0] slv_grp6_p0_w2n_wo_cmd_wmask  ;
  wire    [   2:   0] slv_grp6_p0_w2n_wo_cmd_size   ;
  wire                slv_grp6_p0_w2n_wo_cmd_lock   ;
  wire                slv_grp6_p0_w2n_wo_cmd_excl   ;
  wire    [   7:   0] slv_grp6_p0_w2n_wo_cmd_xlen   ;
  wire    [   1:   0] slv_grp6_p0_w2n_wo_cmd_xburst ;
  wire    [   1:   0] slv_grp6_p0_w2n_wo_cmd_modes  ;
  wire                slv_grp6_p0_w2n_wo_cmd_dmode  ;
  wire    [   2:   0] slv_grp6_p0_w2n_wo_cmd_attri  ;
  wire    [   1:   0] slv_grp6_p0_w2n_wo_cmd_beat   ;
  wire    [   2:   0] slv_grp6_p0_w2n_wo_cmd_usr    ;
  wire                slv_grp6_p0_w2n_wo_rsp_ready  ;
  wire                slv_grp6_p0_w2n_wo_rsp_valid  ;
  wire                slv_grp6_p0_w2n_wo_rsp_err    ;
  wire                slv_grp6_p0_w2n_wo_rsp_excl_ok ;
  wire    [  63:   0] slv_grp6_p0_w2n_wo_rsp_rdata  ;
  wire    [   2:   0] slv_grp6_p0_w2n_wo_rsp_usr    ;
                wire                      slv_grp6_p0_w2n_wo_rsp_last;
   e603_subsys_sgrp6_ficb1ton_bus #(
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (0),
      .ICB_FIFO_CMD_DP        (8),
      .ICB_FIFO_RSP_DP        (8),
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR      (0),
      .O0_BASE_REGION_LSB(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SPLT_FIFO_OUTS_NUM  (8 ),
      .SPLT_FIFO_OUTS_CNT_W(4),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_slv_grp6_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (slv_grp_6_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (slv_grp_6_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (slv_grp_6_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (slv_grp_6_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (slv_grp_6_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp_6_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp_6_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (slv_grp_6_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp_6_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (slv_grp_6_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (slv_grp_6_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp_6_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (slv_grp_6_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp_6_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (slv_grp_6_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp_6_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp_6_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (slv_grp_6_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (slv_grp_6_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (slv_grp_6_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (slv_grp_6_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (slv_grp_6_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp_6_icb_rsp_usr         [   2:   0]),
      .o0_icb_cmd_valid               (slv_grp6_p0_cmd_valid                    ),
  .o0_icb_cmd_ready               (slv_grp6_p0_cmd_ready                    ),
  .o0_icb_cmd_sel                 (slv_grp6_p0_cmd_sel                      ),
  .o0_icb_cmd_read                (slv_grp6_p0_cmd_read                     ),
  .o0_icb_cmd_addr                (slv_grp6_p0_cmd_addr          [  31:   0]),
  .o0_icb_cmd_wdata               (slv_grp6_p0_cmd_wdata         [  63:   0]),
  .o0_icb_cmd_wmask               (slv_grp6_p0_cmd_wmask         [   7:   0]),
  .o0_icb_cmd_size                (slv_grp6_p0_cmd_size          [   2:   0]),
  .o0_icb_cmd_lock                (slv_grp6_p0_cmd_lock                     ),
  .o0_icb_cmd_excl                (slv_grp6_p0_cmd_excl                     ),
  .o0_icb_cmd_xlen                (slv_grp6_p0_cmd_xlen          [   7:   0]),
  .o0_icb_cmd_xburst              (slv_grp6_p0_cmd_xburst        [   1:   0]),
  .o0_icb_cmd_modes               (slv_grp6_p0_cmd_modes         [   1:   0]),
  .o0_icb_cmd_dmode               (slv_grp6_p0_cmd_dmode                    ),
  .o0_icb_cmd_attri               (slv_grp6_p0_cmd_attri         [   2:   0]),
  .o0_icb_cmd_beat                (slv_grp6_p0_cmd_beat          [   1:   0]),
  .o0_icb_cmd_usr                 (slv_grp6_p0_cmd_usr           [   2:   0]),
  .o0_icb_rsp_ready               (slv_grp6_p0_rsp_ready                    ),
  .o0_icb_rsp_valid               (slv_grp6_p0_rsp_valid                    ),
  .o0_icb_rsp_err                 (slv_grp6_p0_rsp_err                      ),
  .o0_icb_rsp_excl_ok             (slv_grp6_p0_rsp_excl_ok                  ),
  .o0_icb_rsp_rdata               (slv_grp6_p0_rsp_rdata         [  63:   0]),
  .o0_icb_rsp_usr                 (slv_grp6_p0_rsp_usr           [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_wconv # (
      .AW    (32),
      .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .ZEROCYC_RSP   (0),
      .FIFO_OUTS_NUM (8),
      .FIFO_CUT_READY(1),
      .X_W(64),
      .Y_W(64 ),
      .CMD_UW (3),
      .RSP_UW (3)
    )u_dummy_slv_icb_icb_wconv(
        .i_icb_cmd_valid                (slv_grp6_p0_cmd_valid                    ),
  .i_icb_cmd_ready                (slv_grp6_p0_cmd_ready                    ),
  .i_icb_cmd_sel                  (slv_grp6_p0_cmd_sel                      ),
  .i_icb_cmd_read                 (slv_grp6_p0_cmd_read                     ),
  .i_icb_cmd_addr                 (slv_grp6_p0_cmd_addr          [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp6_p0_cmd_wdata         [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp6_p0_cmd_wmask         [   7:   0]),
  .i_icb_cmd_size                 (slv_grp6_p0_cmd_size          [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp6_p0_cmd_lock                     ),
  .i_icb_cmd_excl                 (slv_grp6_p0_cmd_excl                     ),
  .i_icb_cmd_xlen                 (slv_grp6_p0_cmd_xlen          [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp6_p0_cmd_xburst        [   1:   0]),
  .i_icb_cmd_modes                (slv_grp6_p0_cmd_modes         [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp6_p0_cmd_dmode                    ),
  .i_icb_cmd_attri                (slv_grp6_p0_cmd_attri         [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp6_p0_cmd_beat          [   1:   0]),
  .i_icb_cmd_usr                  (slv_grp6_p0_cmd_usr           [   2:   0]),
  .i_icb_rsp_ready                (slv_grp6_p0_rsp_ready                    ),
  .i_icb_rsp_valid                (slv_grp6_p0_rsp_valid                    ),
  .i_icb_rsp_err                  (slv_grp6_p0_rsp_err                      ),
  .i_icb_rsp_excl_ok              (slv_grp6_p0_rsp_excl_ok                  ),
  .i_icb_rsp_rdata                (slv_grp6_p0_rsp_rdata         [  63:   0]),
  .i_icb_rsp_usr                  (slv_grp6_p0_rsp_usr           [   2:   0]),
        .o_icb_cmd_valid                (slv_grp6_p0_w2n_cmd_valid                ),
  .o_icb_cmd_ready                (slv_grp6_p0_w2n_cmd_ready                ),
  .o_icb_cmd_sel                  (slv_grp6_p0_w2n_cmd_sel                  ),
  .o_icb_cmd_read                 (slv_grp6_p0_w2n_cmd_read                 ),
  .o_icb_cmd_addr                 (slv_grp6_p0_w2n_cmd_addr      [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp6_p0_w2n_cmd_wdata     [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp6_p0_w2n_cmd_wmask     [   7:   0]),
  .o_icb_cmd_size                 (slv_grp6_p0_w2n_cmd_size      [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp6_p0_w2n_cmd_lock                 ),
  .o_icb_cmd_excl                 (slv_grp6_p0_w2n_cmd_excl                 ),
  .o_icb_cmd_xlen                 (slv_grp6_p0_w2n_cmd_xlen      [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp6_p0_w2n_cmd_xburst    [   1:   0]),
  .o_icb_cmd_modes                (slv_grp6_p0_w2n_cmd_modes     [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp6_p0_w2n_cmd_dmode                ),
  .o_icb_cmd_attri                (slv_grp6_p0_w2n_cmd_attri     [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp6_p0_w2n_cmd_beat      [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp6_p0_w2n_cmd_usr       [   2:   0]),
  .o_icb_rsp_ready                (slv_grp6_p0_w2n_rsp_ready                ),
  .o_icb_rsp_valid                (slv_grp6_p0_w2n_rsp_valid                ),
  .o_icb_rsp_err                  (slv_grp6_p0_w2n_rsp_err                  ),
  .o_icb_rsp_excl_ok              (slv_grp6_p0_w2n_rsp_excl_ok              ),
  .o_icb_rsp_rdata                (slv_grp6_p0_w2n_rsp_rdata     [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp6_p0_w2n_rsp_usr       [   2:   0]),
    .clk  (clk_fab),  
    .rst_n(rst_n)
  );
      assign slv_grp6_p0_w2n_rsp_usr = 3'b0;
      wire dummy_slv_icb_bus_pend_active = 1'b0;
      wire dummy_slv_icb_bus_icb_active;
       e603_subsys_gnrl_ficb_active # (
           .OUTS_CNT_W(4+1)
      )u_dummy_slv_icb__icb_active (
         .icb_active(dummy_slv_icb_bus_icb_active),
            .icb_cmd_valid(slv_grp6_p0_w2n_cmd_valid),
            .icb_cmd_ready(slv_grp6_p0_w2n_cmd_ready),
            .icb_rsp_valid(slv_grp6_p0_w2n_rsp_valid),
            .icb_rsp_ready(slv_grp6_p0_w2n_rsp_ready),
      .clk  (clk_fab),  
      .rst_n(rst_n)
       );
      wire [32-1:0] dummy_slv_icb_cmd_addr_full;
      assign dummy_slv_icb_cmd_addr = dummy_slv_icb_cmd_addr_full[32-1:0];
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(0),
    .O_SUPPORT_RATIO(0),
      .PAYLOAD_NORST(PAYLOAD_NORST),
    .OUTS_CNT_W   (4),
    .AW    (32),
    .DW    (64),
            .CMD_DP    (0),
            .RSP_DP    (0),
            .RSP_BYPBUF(0),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(0),
    .CMD_UW (1),
    .RSP_UW (1)
  )u_dummy_slv_icb_icb_buffer(
    .i_clk_en (1'b1),
    .o_clk_en (1'b1),
    .icb_buffer_active   (),
             .i_icb_cmd_usr(1'b0),
             .i_icb_rsp_usr(),
      .i_icb_cmd_valid                (slv_grp6_p0_w2n_cmd_valid                ),
  .i_icb_cmd_ready                (slv_grp6_p0_w2n_cmd_ready                ),
  .i_icb_cmd_sel                  (slv_grp6_p0_w2n_cmd_sel                  ),
  .i_icb_cmd_read                 (slv_grp6_p0_w2n_cmd_read                 ),
  .i_icb_cmd_addr                 (slv_grp6_p0_w2n_cmd_addr      [  31:   0]),
  .i_icb_cmd_wdata                (slv_grp6_p0_w2n_cmd_wdata     [  63:   0]),
  .i_icb_cmd_wmask                (slv_grp6_p0_w2n_cmd_wmask     [   7:   0]),
  .i_icb_cmd_size                 (slv_grp6_p0_w2n_cmd_size      [   2:   0]),
  .i_icb_cmd_lock                 (slv_grp6_p0_w2n_cmd_lock                 ),
  .i_icb_cmd_excl                 (slv_grp6_p0_w2n_cmd_excl                 ),
  .i_icb_cmd_xlen                 (slv_grp6_p0_w2n_cmd_xlen      [   7:   0]),
  .i_icb_cmd_xburst               (slv_grp6_p0_w2n_cmd_xburst    [   1:   0]),
  .i_icb_cmd_modes                (slv_grp6_p0_w2n_cmd_modes     [   1:   0]),
  .i_icb_cmd_dmode                (slv_grp6_p0_w2n_cmd_dmode                ),
  .i_icb_cmd_attri                (slv_grp6_p0_w2n_cmd_attri     [   2:   0]),
  .i_icb_cmd_beat                 (slv_grp6_p0_w2n_cmd_beat      [   1:   0]),
  .i_icb_rsp_ready                (slv_grp6_p0_w2n_rsp_ready                ),
  .i_icb_rsp_valid                (slv_grp6_p0_w2n_rsp_valid                ),
  .i_icb_rsp_err                  (slv_grp6_p0_w2n_rsp_err                  ),
  .i_icb_rsp_excl_ok              (slv_grp6_p0_w2n_rsp_excl_ok              ),
  .i_icb_rsp_rdata                (slv_grp6_p0_w2n_rsp_rdata     [  63:   0]),
      .o_icb_cmd_valid                (dummy_slv_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (dummy_slv_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (dummy_slv_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (dummy_slv_icb_cmd_read                   ),
  .o_icb_cmd_wdata                (dummy_slv_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (dummy_slv_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (dummy_slv_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (dummy_slv_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (dummy_slv_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (dummy_slv_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (dummy_slv_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (dummy_slv_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (dummy_slv_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (dummy_slv_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (dummy_slv_icb_cmd_beat        [   1:   0]),
  .o_icb_rsp_ready                (dummy_slv_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (dummy_slv_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (dummy_slv_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (dummy_slv_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (dummy_slv_icb_rsp_rdata       [  63:   0]),
            .o_icb_cmd_usr(),
            .o_icb_rsp_usr(1'b0),
      .o_icb_cmd_addr(dummy_slv_icb_cmd_addr_full),
      .clk  (clk_fab),  
      .rst_n(rst_n)
  );
              wire                xbar_mg0_ro_to_sg0_cmd_valid  ;
  wire                xbar_mg0_ro_to_sg0_cmd_ready  ;
  wire                xbar_mg0_ro_to_sg0_cmd_sel    ;
  wire                xbar_mg0_ro_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg0_ro_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_ro_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_ro_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg0_cmd_size   ;
  wire                xbar_mg0_ro_to_sg0_cmd_lock   ;
  wire                xbar_mg0_ro_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_ro_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_ro_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_ro_to_sg0_cmd_modes  ;
  wire                xbar_mg0_ro_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_ro_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_ro_to_sg0_cmd_usr    ;
  wire                xbar_mg0_ro_to_sg0_rsp_ready  ;
  wire                xbar_mg0_ro_to_sg0_rsp_valid  ;
  wire                xbar_mg0_ro_to_sg0_rsp_err    ;
  wire                xbar_mg0_ro_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_ro_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg0_rsp_usr    ;
              wire                xbar_mg0_wo_to_sg0_cmd_valid  ;
  wire                xbar_mg0_wo_to_sg0_cmd_ready  ;
  wire                xbar_mg0_wo_to_sg0_cmd_sel    ;
  wire                xbar_mg0_wo_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg0_wo_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_wo_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_wo_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg0_cmd_size   ;
  wire                xbar_mg0_wo_to_sg0_cmd_lock   ;
  wire                xbar_mg0_wo_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_wo_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_wo_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_wo_to_sg0_cmd_modes  ;
  wire                xbar_mg0_wo_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_wo_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_wo_to_sg0_cmd_usr    ;
  wire                xbar_mg0_wo_to_sg0_rsp_ready  ;
  wire                xbar_mg0_wo_to_sg0_rsp_valid  ;
  wire                xbar_mg0_wo_to_sg0_rsp_err    ;
  wire                xbar_mg0_wo_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_wo_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg0_rsp_usr    ;
              wire                xbar_mg0_ro_to_sg1_cmd_valid  ;
  wire                xbar_mg0_ro_to_sg1_cmd_ready  ;
  wire                xbar_mg0_ro_to_sg1_cmd_sel    ;
  wire                xbar_mg0_ro_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg0_ro_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_ro_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_ro_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg1_cmd_size   ;
  wire                xbar_mg0_ro_to_sg1_cmd_lock   ;
  wire                xbar_mg0_ro_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_ro_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_ro_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_ro_to_sg1_cmd_modes  ;
  wire                xbar_mg0_ro_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_ro_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_ro_to_sg1_cmd_usr    ;
  wire                xbar_mg0_ro_to_sg1_rsp_ready  ;
  wire                xbar_mg0_ro_to_sg1_rsp_valid  ;
  wire                xbar_mg0_ro_to_sg1_rsp_err    ;
  wire                xbar_mg0_ro_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_ro_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg1_rsp_usr    ;
              wire                xbar_mg0_wo_to_sg1_cmd_valid  ;
  wire                xbar_mg0_wo_to_sg1_cmd_ready  ;
  wire                xbar_mg0_wo_to_sg1_cmd_sel    ;
  wire                xbar_mg0_wo_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg0_wo_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_wo_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_wo_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg1_cmd_size   ;
  wire                xbar_mg0_wo_to_sg1_cmd_lock   ;
  wire                xbar_mg0_wo_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_wo_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_wo_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_wo_to_sg1_cmd_modes  ;
  wire                xbar_mg0_wo_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_wo_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_wo_to_sg1_cmd_usr    ;
  wire                xbar_mg0_wo_to_sg1_rsp_ready  ;
  wire                xbar_mg0_wo_to_sg1_rsp_valid  ;
  wire                xbar_mg0_wo_to_sg1_rsp_err    ;
  wire                xbar_mg0_wo_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_wo_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg1_rsp_usr    ;
              wire                xbar_mg0_ro_to_sg2_cmd_valid  ;
  wire                xbar_mg0_ro_to_sg2_cmd_ready  ;
  wire                xbar_mg0_ro_to_sg2_cmd_sel    ;
  wire                xbar_mg0_ro_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg0_ro_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_ro_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_ro_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg2_cmd_size   ;
  wire                xbar_mg0_ro_to_sg2_cmd_lock   ;
  wire                xbar_mg0_ro_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_ro_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_ro_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_ro_to_sg2_cmd_modes  ;
  wire                xbar_mg0_ro_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_ro_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_ro_to_sg2_cmd_usr    ;
  wire                xbar_mg0_ro_to_sg2_rsp_ready  ;
  wire                xbar_mg0_ro_to_sg2_rsp_valid  ;
  wire                xbar_mg0_ro_to_sg2_rsp_err    ;
  wire                xbar_mg0_ro_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_ro_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg2_rsp_usr    ;
              wire                xbar_mg0_wo_to_sg2_cmd_valid  ;
  wire                xbar_mg0_wo_to_sg2_cmd_ready  ;
  wire                xbar_mg0_wo_to_sg2_cmd_sel    ;
  wire                xbar_mg0_wo_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg0_wo_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_wo_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_wo_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg2_cmd_size   ;
  wire                xbar_mg0_wo_to_sg2_cmd_lock   ;
  wire                xbar_mg0_wo_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_wo_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_wo_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_wo_to_sg2_cmd_modes  ;
  wire                xbar_mg0_wo_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_wo_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_wo_to_sg2_cmd_usr    ;
  wire                xbar_mg0_wo_to_sg2_rsp_ready  ;
  wire                xbar_mg0_wo_to_sg2_rsp_valid  ;
  wire                xbar_mg0_wo_to_sg2_rsp_err    ;
  wire                xbar_mg0_wo_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_wo_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg2_rsp_usr    ;
              wire                xbar_mg0_ro_to_sg3_cmd_valid  ;
  wire                xbar_mg0_ro_to_sg3_cmd_ready  ;
  wire                xbar_mg0_ro_to_sg3_cmd_sel    ;
  wire                xbar_mg0_ro_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg0_ro_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_ro_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_ro_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg3_cmd_size   ;
  wire                xbar_mg0_ro_to_sg3_cmd_lock   ;
  wire                xbar_mg0_ro_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_ro_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_ro_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_ro_to_sg3_cmd_modes  ;
  wire                xbar_mg0_ro_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_ro_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_ro_to_sg3_cmd_usr    ;
  wire                xbar_mg0_ro_to_sg3_rsp_ready  ;
  wire                xbar_mg0_ro_to_sg3_rsp_valid  ;
  wire                xbar_mg0_ro_to_sg3_rsp_err    ;
  wire                xbar_mg0_ro_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_ro_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg3_rsp_usr    ;
              wire                xbar_mg0_wo_to_sg3_cmd_valid  ;
  wire                xbar_mg0_wo_to_sg3_cmd_ready  ;
  wire                xbar_mg0_wo_to_sg3_cmd_sel    ;
  wire                xbar_mg0_wo_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg0_wo_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_wo_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_wo_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg3_cmd_size   ;
  wire                xbar_mg0_wo_to_sg3_cmd_lock   ;
  wire                xbar_mg0_wo_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_wo_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_wo_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_wo_to_sg3_cmd_modes  ;
  wire                xbar_mg0_wo_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_wo_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_wo_to_sg3_cmd_usr    ;
  wire                xbar_mg0_wo_to_sg3_rsp_ready  ;
  wire                xbar_mg0_wo_to_sg3_rsp_valid  ;
  wire                xbar_mg0_wo_to_sg3_rsp_err    ;
  wire                xbar_mg0_wo_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_wo_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg3_rsp_usr    ;
              wire                xbar_mg0_ro_to_sg4_cmd_valid  ;
  wire                xbar_mg0_ro_to_sg4_cmd_ready  ;
  wire                xbar_mg0_ro_to_sg4_cmd_sel    ;
  wire                xbar_mg0_ro_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg0_ro_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_ro_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_ro_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg4_cmd_size   ;
  wire                xbar_mg0_ro_to_sg4_cmd_lock   ;
  wire                xbar_mg0_ro_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_ro_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_ro_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_ro_to_sg4_cmd_modes  ;
  wire                xbar_mg0_ro_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_ro_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_ro_to_sg4_cmd_usr    ;
  wire                xbar_mg0_ro_to_sg4_rsp_ready  ;
  wire                xbar_mg0_ro_to_sg4_rsp_valid  ;
  wire                xbar_mg0_ro_to_sg4_rsp_err    ;
  wire                xbar_mg0_ro_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_ro_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg4_rsp_usr    ;
              wire                xbar_mg0_wo_to_sg4_cmd_valid  ;
  wire                xbar_mg0_wo_to_sg4_cmd_ready  ;
  wire                xbar_mg0_wo_to_sg4_cmd_sel    ;
  wire                xbar_mg0_wo_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg0_wo_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_wo_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_wo_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg4_cmd_size   ;
  wire                xbar_mg0_wo_to_sg4_cmd_lock   ;
  wire                xbar_mg0_wo_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_wo_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_wo_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_wo_to_sg4_cmd_modes  ;
  wire                xbar_mg0_wo_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_wo_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_wo_to_sg4_cmd_usr    ;
  wire                xbar_mg0_wo_to_sg4_rsp_ready  ;
  wire                xbar_mg0_wo_to_sg4_rsp_valid  ;
  wire                xbar_mg0_wo_to_sg4_rsp_err    ;
  wire                xbar_mg0_wo_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_wo_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg4_rsp_usr    ;
              wire                xbar_mg0_ro_to_sg5_cmd_valid  ;
  wire                xbar_mg0_ro_to_sg5_cmd_ready  ;
  wire                xbar_mg0_ro_to_sg5_cmd_sel    ;
  wire                xbar_mg0_ro_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg0_ro_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_ro_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_ro_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg5_cmd_size   ;
  wire                xbar_mg0_ro_to_sg5_cmd_lock   ;
  wire                xbar_mg0_ro_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_ro_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_ro_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_ro_to_sg5_cmd_modes  ;
  wire                xbar_mg0_ro_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_ro_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_ro_to_sg5_cmd_usr    ;
  wire                xbar_mg0_ro_to_sg5_rsp_ready  ;
  wire                xbar_mg0_ro_to_sg5_rsp_valid  ;
  wire                xbar_mg0_ro_to_sg5_rsp_err    ;
  wire                xbar_mg0_ro_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_ro_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg5_rsp_usr    ;
              wire                xbar_mg0_wo_to_sg5_cmd_valid  ;
  wire                xbar_mg0_wo_to_sg5_cmd_ready  ;
  wire                xbar_mg0_wo_to_sg5_cmd_sel    ;
  wire                xbar_mg0_wo_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg0_wo_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_wo_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_wo_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg5_cmd_size   ;
  wire                xbar_mg0_wo_to_sg5_cmd_lock   ;
  wire                xbar_mg0_wo_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_wo_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_wo_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_wo_to_sg5_cmd_modes  ;
  wire                xbar_mg0_wo_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_wo_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_wo_to_sg5_cmd_usr    ;
  wire                xbar_mg0_wo_to_sg5_rsp_ready  ;
  wire                xbar_mg0_wo_to_sg5_rsp_valid  ;
  wire                xbar_mg0_wo_to_sg5_rsp_err    ;
  wire                xbar_mg0_wo_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_wo_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg5_rsp_usr    ;
              wire                xbar_mg0_ro_to_sg6_cmd_valid  ;
  wire                xbar_mg0_ro_to_sg6_cmd_ready  ;
  wire                xbar_mg0_ro_to_sg6_cmd_sel    ;
  wire                xbar_mg0_ro_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg0_ro_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_ro_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_ro_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg6_cmd_size   ;
  wire                xbar_mg0_ro_to_sg6_cmd_lock   ;
  wire                xbar_mg0_ro_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_ro_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_ro_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_ro_to_sg6_cmd_modes  ;
  wire                xbar_mg0_ro_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_ro_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_ro_to_sg6_cmd_usr    ;
  wire                xbar_mg0_ro_to_sg6_rsp_ready  ;
  wire                xbar_mg0_ro_to_sg6_rsp_valid  ;
  wire                xbar_mg0_ro_to_sg6_rsp_err    ;
  wire                xbar_mg0_ro_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_ro_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_ro_to_sg6_rsp_usr    ;
              wire                xbar_mg0_wo_to_sg6_cmd_valid  ;
  wire                xbar_mg0_wo_to_sg6_cmd_ready  ;
  wire                xbar_mg0_wo_to_sg6_cmd_sel    ;
  wire                xbar_mg0_wo_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg0_wo_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg0_wo_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg0_wo_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg6_cmd_size   ;
  wire                xbar_mg0_wo_to_sg6_cmd_lock   ;
  wire                xbar_mg0_wo_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg0_wo_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg0_wo_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg0_wo_to_sg6_cmd_modes  ;
  wire                xbar_mg0_wo_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg0_wo_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg0_wo_to_sg6_cmd_usr    ;
  wire                xbar_mg0_wo_to_sg6_rsp_ready  ;
  wire                xbar_mg0_wo_to_sg6_rsp_valid  ;
  wire                xbar_mg0_wo_to_sg6_rsp_err    ;
  wire                xbar_mg0_wo_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg0_wo_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg0_wo_to_sg6_rsp_usr    ;
              wire                xbar_mg1_ro_to_sg0_cmd_valid  ;
  wire                xbar_mg1_ro_to_sg0_cmd_ready  ;
  wire                xbar_mg1_ro_to_sg0_cmd_sel    ;
  wire                xbar_mg1_ro_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg1_ro_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg1_ro_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg1_ro_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg0_cmd_size   ;
  wire                xbar_mg1_ro_to_sg0_cmd_lock   ;
  wire                xbar_mg1_ro_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg1_ro_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg1_ro_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg1_ro_to_sg0_cmd_modes  ;
  wire                xbar_mg1_ro_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg1_ro_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg1_ro_to_sg0_cmd_usr    ;
  wire                xbar_mg1_ro_to_sg0_rsp_ready  ;
  wire                xbar_mg1_ro_to_sg0_rsp_valid  ;
  wire                xbar_mg1_ro_to_sg0_rsp_err    ;
  wire                xbar_mg1_ro_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg1_ro_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg0_rsp_usr    ;
              wire                xbar_mg1_ro_to_sg1_cmd_valid  ;
  wire                xbar_mg1_ro_to_sg1_cmd_ready  ;
  wire                xbar_mg1_ro_to_sg1_cmd_sel    ;
  wire                xbar_mg1_ro_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg1_ro_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg1_ro_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg1_ro_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg1_cmd_size   ;
  wire                xbar_mg1_ro_to_sg1_cmd_lock   ;
  wire                xbar_mg1_ro_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg1_ro_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg1_ro_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg1_ro_to_sg1_cmd_modes  ;
  wire                xbar_mg1_ro_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg1_ro_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg1_ro_to_sg1_cmd_usr    ;
  wire                xbar_mg1_ro_to_sg1_rsp_ready  ;
  wire                xbar_mg1_ro_to_sg1_rsp_valid  ;
  wire                xbar_mg1_ro_to_sg1_rsp_err    ;
  wire                xbar_mg1_ro_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg1_ro_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg1_rsp_usr    ;
              wire                xbar_mg1_ro_to_sg2_cmd_valid  ;
  wire                xbar_mg1_ro_to_sg2_cmd_ready  ;
  wire                xbar_mg1_ro_to_sg2_cmd_sel    ;
  wire                xbar_mg1_ro_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg1_ro_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg1_ro_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg1_ro_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg2_cmd_size   ;
  wire                xbar_mg1_ro_to_sg2_cmd_lock   ;
  wire                xbar_mg1_ro_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg1_ro_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg1_ro_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg1_ro_to_sg2_cmd_modes  ;
  wire                xbar_mg1_ro_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg1_ro_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg1_ro_to_sg2_cmd_usr    ;
  wire                xbar_mg1_ro_to_sg2_rsp_ready  ;
  wire                xbar_mg1_ro_to_sg2_rsp_valid  ;
  wire                xbar_mg1_ro_to_sg2_rsp_err    ;
  wire                xbar_mg1_ro_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg1_ro_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg2_rsp_usr    ;
              wire                xbar_mg1_ro_to_sg3_cmd_valid  ;
  wire                xbar_mg1_ro_to_sg3_cmd_ready  ;
  wire                xbar_mg1_ro_to_sg3_cmd_sel    ;
  wire                xbar_mg1_ro_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg1_ro_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg1_ro_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg1_ro_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg3_cmd_size   ;
  wire                xbar_mg1_ro_to_sg3_cmd_lock   ;
  wire                xbar_mg1_ro_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg1_ro_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg1_ro_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg1_ro_to_sg3_cmd_modes  ;
  wire                xbar_mg1_ro_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg1_ro_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg1_ro_to_sg3_cmd_usr    ;
  wire                xbar_mg1_ro_to_sg3_rsp_ready  ;
  wire                xbar_mg1_ro_to_sg3_rsp_valid  ;
  wire                xbar_mg1_ro_to_sg3_rsp_err    ;
  wire                xbar_mg1_ro_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg1_ro_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg3_rsp_usr    ;
              wire                xbar_mg1_ro_to_sg4_cmd_valid  ;
  wire                xbar_mg1_ro_to_sg4_cmd_ready  ;
  wire                xbar_mg1_ro_to_sg4_cmd_sel    ;
  wire                xbar_mg1_ro_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg1_ro_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg1_ro_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg1_ro_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg4_cmd_size   ;
  wire                xbar_mg1_ro_to_sg4_cmd_lock   ;
  wire                xbar_mg1_ro_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg1_ro_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg1_ro_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg1_ro_to_sg4_cmd_modes  ;
  wire                xbar_mg1_ro_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg1_ro_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg1_ro_to_sg4_cmd_usr    ;
  wire                xbar_mg1_ro_to_sg4_rsp_ready  ;
  wire                xbar_mg1_ro_to_sg4_rsp_valid  ;
  wire                xbar_mg1_ro_to_sg4_rsp_err    ;
  wire                xbar_mg1_ro_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg1_ro_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg4_rsp_usr    ;
              wire                xbar_mg1_ro_to_sg5_cmd_valid  ;
  wire                xbar_mg1_ro_to_sg5_cmd_ready  ;
  wire                xbar_mg1_ro_to_sg5_cmd_sel    ;
  wire                xbar_mg1_ro_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg1_ro_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg1_ro_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg1_ro_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg5_cmd_size   ;
  wire                xbar_mg1_ro_to_sg5_cmd_lock   ;
  wire                xbar_mg1_ro_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg1_ro_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg1_ro_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg1_ro_to_sg5_cmd_modes  ;
  wire                xbar_mg1_ro_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg1_ro_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg1_ro_to_sg5_cmd_usr    ;
  wire                xbar_mg1_ro_to_sg5_rsp_ready  ;
  wire                xbar_mg1_ro_to_sg5_rsp_valid  ;
  wire                xbar_mg1_ro_to_sg5_rsp_err    ;
  wire                xbar_mg1_ro_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg1_ro_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg5_rsp_usr    ;
              wire                xbar_mg1_ro_to_sg6_cmd_valid  ;
  wire                xbar_mg1_ro_to_sg6_cmd_ready  ;
  wire                xbar_mg1_ro_to_sg6_cmd_sel    ;
  wire                xbar_mg1_ro_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg1_ro_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg1_ro_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg1_ro_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg6_cmd_size   ;
  wire                xbar_mg1_ro_to_sg6_cmd_lock   ;
  wire                xbar_mg1_ro_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg1_ro_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg1_ro_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg1_ro_to_sg6_cmd_modes  ;
  wire                xbar_mg1_ro_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg1_ro_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg1_ro_to_sg6_cmd_usr    ;
  wire                xbar_mg1_ro_to_sg6_rsp_ready  ;
  wire                xbar_mg1_ro_to_sg6_rsp_valid  ;
  wire                xbar_mg1_ro_to_sg6_rsp_err    ;
  wire                xbar_mg1_ro_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg1_ro_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg1_ro_to_sg6_rsp_usr    ;
              wire                xbar_mg2_wo_to_sg0_cmd_valid  ;
  wire                xbar_mg2_wo_to_sg0_cmd_ready  ;
  wire                xbar_mg2_wo_to_sg0_cmd_sel    ;
  wire                xbar_mg2_wo_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg2_wo_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg2_wo_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg2_wo_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg0_cmd_size   ;
  wire                xbar_mg2_wo_to_sg0_cmd_lock   ;
  wire                xbar_mg2_wo_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg2_wo_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg2_wo_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg2_wo_to_sg0_cmd_modes  ;
  wire                xbar_mg2_wo_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg2_wo_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg2_wo_to_sg0_cmd_usr    ;
  wire                xbar_mg2_wo_to_sg0_rsp_ready  ;
  wire                xbar_mg2_wo_to_sg0_rsp_valid  ;
  wire                xbar_mg2_wo_to_sg0_rsp_err    ;
  wire                xbar_mg2_wo_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg2_wo_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg0_rsp_usr    ;
              wire                xbar_mg2_wo_to_sg1_cmd_valid  ;
  wire                xbar_mg2_wo_to_sg1_cmd_ready  ;
  wire                xbar_mg2_wo_to_sg1_cmd_sel    ;
  wire                xbar_mg2_wo_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg2_wo_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg2_wo_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg2_wo_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg1_cmd_size   ;
  wire                xbar_mg2_wo_to_sg1_cmd_lock   ;
  wire                xbar_mg2_wo_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg2_wo_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg2_wo_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg2_wo_to_sg1_cmd_modes  ;
  wire                xbar_mg2_wo_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg2_wo_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg2_wo_to_sg1_cmd_usr    ;
  wire                xbar_mg2_wo_to_sg1_rsp_ready  ;
  wire                xbar_mg2_wo_to_sg1_rsp_valid  ;
  wire                xbar_mg2_wo_to_sg1_rsp_err    ;
  wire                xbar_mg2_wo_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg2_wo_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg1_rsp_usr    ;
              wire                xbar_mg2_wo_to_sg2_cmd_valid  ;
  wire                xbar_mg2_wo_to_sg2_cmd_ready  ;
  wire                xbar_mg2_wo_to_sg2_cmd_sel    ;
  wire                xbar_mg2_wo_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg2_wo_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg2_wo_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg2_wo_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg2_cmd_size   ;
  wire                xbar_mg2_wo_to_sg2_cmd_lock   ;
  wire                xbar_mg2_wo_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg2_wo_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg2_wo_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg2_wo_to_sg2_cmd_modes  ;
  wire                xbar_mg2_wo_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg2_wo_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg2_wo_to_sg2_cmd_usr    ;
  wire                xbar_mg2_wo_to_sg2_rsp_ready  ;
  wire                xbar_mg2_wo_to_sg2_rsp_valid  ;
  wire                xbar_mg2_wo_to_sg2_rsp_err    ;
  wire                xbar_mg2_wo_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg2_wo_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg2_rsp_usr    ;
              wire                xbar_mg2_wo_to_sg3_cmd_valid  ;
  wire                xbar_mg2_wo_to_sg3_cmd_ready  ;
  wire                xbar_mg2_wo_to_sg3_cmd_sel    ;
  wire                xbar_mg2_wo_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg2_wo_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg2_wo_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg2_wo_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg3_cmd_size   ;
  wire                xbar_mg2_wo_to_sg3_cmd_lock   ;
  wire                xbar_mg2_wo_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg2_wo_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg2_wo_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg2_wo_to_sg3_cmd_modes  ;
  wire                xbar_mg2_wo_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg2_wo_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg2_wo_to_sg3_cmd_usr    ;
  wire                xbar_mg2_wo_to_sg3_rsp_ready  ;
  wire                xbar_mg2_wo_to_sg3_rsp_valid  ;
  wire                xbar_mg2_wo_to_sg3_rsp_err    ;
  wire                xbar_mg2_wo_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg2_wo_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg3_rsp_usr    ;
              wire                xbar_mg2_wo_to_sg4_cmd_valid  ;
  wire                xbar_mg2_wo_to_sg4_cmd_ready  ;
  wire                xbar_mg2_wo_to_sg4_cmd_sel    ;
  wire                xbar_mg2_wo_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg2_wo_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg2_wo_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg2_wo_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg4_cmd_size   ;
  wire                xbar_mg2_wo_to_sg4_cmd_lock   ;
  wire                xbar_mg2_wo_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg2_wo_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg2_wo_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg2_wo_to_sg4_cmd_modes  ;
  wire                xbar_mg2_wo_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg2_wo_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg2_wo_to_sg4_cmd_usr    ;
  wire                xbar_mg2_wo_to_sg4_rsp_ready  ;
  wire                xbar_mg2_wo_to_sg4_rsp_valid  ;
  wire                xbar_mg2_wo_to_sg4_rsp_err    ;
  wire                xbar_mg2_wo_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg2_wo_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg4_rsp_usr    ;
              wire                xbar_mg2_wo_to_sg5_cmd_valid  ;
  wire                xbar_mg2_wo_to_sg5_cmd_ready  ;
  wire                xbar_mg2_wo_to_sg5_cmd_sel    ;
  wire                xbar_mg2_wo_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg2_wo_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg2_wo_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg2_wo_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg5_cmd_size   ;
  wire                xbar_mg2_wo_to_sg5_cmd_lock   ;
  wire                xbar_mg2_wo_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg2_wo_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg2_wo_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg2_wo_to_sg5_cmd_modes  ;
  wire                xbar_mg2_wo_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg2_wo_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg2_wo_to_sg5_cmd_usr    ;
  wire                xbar_mg2_wo_to_sg5_rsp_ready  ;
  wire                xbar_mg2_wo_to_sg5_rsp_valid  ;
  wire                xbar_mg2_wo_to_sg5_rsp_err    ;
  wire                xbar_mg2_wo_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg2_wo_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg5_rsp_usr    ;
              wire                xbar_mg2_wo_to_sg6_cmd_valid  ;
  wire                xbar_mg2_wo_to_sg6_cmd_ready  ;
  wire                xbar_mg2_wo_to_sg6_cmd_sel    ;
  wire                xbar_mg2_wo_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg2_wo_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg2_wo_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg2_wo_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg6_cmd_size   ;
  wire                xbar_mg2_wo_to_sg6_cmd_lock   ;
  wire                xbar_mg2_wo_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg2_wo_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg2_wo_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg2_wo_to_sg6_cmd_modes  ;
  wire                xbar_mg2_wo_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg2_wo_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg2_wo_to_sg6_cmd_usr    ;
  wire                xbar_mg2_wo_to_sg6_rsp_ready  ;
  wire                xbar_mg2_wo_to_sg6_rsp_valid  ;
  wire                xbar_mg2_wo_to_sg6_rsp_err    ;
  wire                xbar_mg2_wo_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg2_wo_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg2_wo_to_sg6_rsp_usr    ;
              wire                xbar_mg3_ro_to_sg0_cmd_valid  ;
  wire                xbar_mg3_ro_to_sg0_cmd_ready  ;
  wire                xbar_mg3_ro_to_sg0_cmd_sel    ;
  wire                xbar_mg3_ro_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg3_ro_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_ro_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_ro_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg0_cmd_size   ;
  wire                xbar_mg3_ro_to_sg0_cmd_lock   ;
  wire                xbar_mg3_ro_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_ro_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_ro_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_ro_to_sg0_cmd_modes  ;
  wire                xbar_mg3_ro_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_ro_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_ro_to_sg0_cmd_usr    ;
  wire                xbar_mg3_ro_to_sg0_rsp_ready  ;
  wire                xbar_mg3_ro_to_sg0_rsp_valid  ;
  wire                xbar_mg3_ro_to_sg0_rsp_err    ;
  wire                xbar_mg3_ro_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_ro_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg0_rsp_usr    ;
              wire                xbar_mg3_wo_to_sg0_cmd_valid  ;
  wire                xbar_mg3_wo_to_sg0_cmd_ready  ;
  wire                xbar_mg3_wo_to_sg0_cmd_sel    ;
  wire                xbar_mg3_wo_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg3_wo_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_wo_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_wo_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg0_cmd_size   ;
  wire                xbar_mg3_wo_to_sg0_cmd_lock   ;
  wire                xbar_mg3_wo_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_wo_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_wo_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_wo_to_sg0_cmd_modes  ;
  wire                xbar_mg3_wo_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_wo_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_wo_to_sg0_cmd_usr    ;
  wire                xbar_mg3_wo_to_sg0_rsp_ready  ;
  wire                xbar_mg3_wo_to_sg0_rsp_valid  ;
  wire                xbar_mg3_wo_to_sg0_rsp_err    ;
  wire                xbar_mg3_wo_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_wo_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg0_rsp_usr    ;
              wire                xbar_mg3_ro_to_sg1_cmd_valid  ;
  wire                xbar_mg3_ro_to_sg1_cmd_ready  ;
  wire                xbar_mg3_ro_to_sg1_cmd_sel    ;
  wire                xbar_mg3_ro_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg3_ro_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_ro_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_ro_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg1_cmd_size   ;
  wire                xbar_mg3_ro_to_sg1_cmd_lock   ;
  wire                xbar_mg3_ro_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_ro_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_ro_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_ro_to_sg1_cmd_modes  ;
  wire                xbar_mg3_ro_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_ro_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_ro_to_sg1_cmd_usr    ;
  wire                xbar_mg3_ro_to_sg1_rsp_ready  ;
  wire                xbar_mg3_ro_to_sg1_rsp_valid  ;
  wire                xbar_mg3_ro_to_sg1_rsp_err    ;
  wire                xbar_mg3_ro_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_ro_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg1_rsp_usr    ;
              wire                xbar_mg3_wo_to_sg1_cmd_valid  ;
  wire                xbar_mg3_wo_to_sg1_cmd_ready  ;
  wire                xbar_mg3_wo_to_sg1_cmd_sel    ;
  wire                xbar_mg3_wo_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg3_wo_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_wo_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_wo_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg1_cmd_size   ;
  wire                xbar_mg3_wo_to_sg1_cmd_lock   ;
  wire                xbar_mg3_wo_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_wo_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_wo_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_wo_to_sg1_cmd_modes  ;
  wire                xbar_mg3_wo_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_wo_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_wo_to_sg1_cmd_usr    ;
  wire                xbar_mg3_wo_to_sg1_rsp_ready  ;
  wire                xbar_mg3_wo_to_sg1_rsp_valid  ;
  wire                xbar_mg3_wo_to_sg1_rsp_err    ;
  wire                xbar_mg3_wo_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_wo_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg1_rsp_usr    ;
              wire                xbar_mg3_ro_to_sg2_cmd_valid  ;
  wire                xbar_mg3_ro_to_sg2_cmd_ready  ;
  wire                xbar_mg3_ro_to_sg2_cmd_sel    ;
  wire                xbar_mg3_ro_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg3_ro_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_ro_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_ro_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg2_cmd_size   ;
  wire                xbar_mg3_ro_to_sg2_cmd_lock   ;
  wire                xbar_mg3_ro_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_ro_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_ro_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_ro_to_sg2_cmd_modes  ;
  wire                xbar_mg3_ro_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_ro_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_ro_to_sg2_cmd_usr    ;
  wire                xbar_mg3_ro_to_sg2_rsp_ready  ;
  wire                xbar_mg3_ro_to_sg2_rsp_valid  ;
  wire                xbar_mg3_ro_to_sg2_rsp_err    ;
  wire                xbar_mg3_ro_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_ro_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg2_rsp_usr    ;
              wire                xbar_mg3_wo_to_sg2_cmd_valid  ;
  wire                xbar_mg3_wo_to_sg2_cmd_ready  ;
  wire                xbar_mg3_wo_to_sg2_cmd_sel    ;
  wire                xbar_mg3_wo_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg3_wo_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_wo_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_wo_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg2_cmd_size   ;
  wire                xbar_mg3_wo_to_sg2_cmd_lock   ;
  wire                xbar_mg3_wo_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_wo_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_wo_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_wo_to_sg2_cmd_modes  ;
  wire                xbar_mg3_wo_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_wo_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_wo_to_sg2_cmd_usr    ;
  wire                xbar_mg3_wo_to_sg2_rsp_ready  ;
  wire                xbar_mg3_wo_to_sg2_rsp_valid  ;
  wire                xbar_mg3_wo_to_sg2_rsp_err    ;
  wire                xbar_mg3_wo_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_wo_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg2_rsp_usr    ;
              wire                xbar_mg3_ro_to_sg3_cmd_valid  ;
  wire                xbar_mg3_ro_to_sg3_cmd_ready  ;
  wire                xbar_mg3_ro_to_sg3_cmd_sel    ;
  wire                xbar_mg3_ro_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg3_ro_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_ro_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_ro_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg3_cmd_size   ;
  wire                xbar_mg3_ro_to_sg3_cmd_lock   ;
  wire                xbar_mg3_ro_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_ro_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_ro_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_ro_to_sg3_cmd_modes  ;
  wire                xbar_mg3_ro_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_ro_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_ro_to_sg3_cmd_usr    ;
  wire                xbar_mg3_ro_to_sg3_rsp_ready  ;
  wire                xbar_mg3_ro_to_sg3_rsp_valid  ;
  wire                xbar_mg3_ro_to_sg3_rsp_err    ;
  wire                xbar_mg3_ro_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_ro_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg3_rsp_usr    ;
              wire                xbar_mg3_wo_to_sg3_cmd_valid  ;
  wire                xbar_mg3_wo_to_sg3_cmd_ready  ;
  wire                xbar_mg3_wo_to_sg3_cmd_sel    ;
  wire                xbar_mg3_wo_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg3_wo_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_wo_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_wo_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg3_cmd_size   ;
  wire                xbar_mg3_wo_to_sg3_cmd_lock   ;
  wire                xbar_mg3_wo_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_wo_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_wo_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_wo_to_sg3_cmd_modes  ;
  wire                xbar_mg3_wo_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_wo_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_wo_to_sg3_cmd_usr    ;
  wire                xbar_mg3_wo_to_sg3_rsp_ready  ;
  wire                xbar_mg3_wo_to_sg3_rsp_valid  ;
  wire                xbar_mg3_wo_to_sg3_rsp_err    ;
  wire                xbar_mg3_wo_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_wo_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg3_rsp_usr    ;
              wire                xbar_mg3_ro_to_sg4_cmd_valid  ;
  wire                xbar_mg3_ro_to_sg4_cmd_ready  ;
  wire                xbar_mg3_ro_to_sg4_cmd_sel    ;
  wire                xbar_mg3_ro_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg3_ro_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_ro_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_ro_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg4_cmd_size   ;
  wire                xbar_mg3_ro_to_sg4_cmd_lock   ;
  wire                xbar_mg3_ro_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_ro_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_ro_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_ro_to_sg4_cmd_modes  ;
  wire                xbar_mg3_ro_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_ro_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_ro_to_sg4_cmd_usr    ;
  wire                xbar_mg3_ro_to_sg4_rsp_ready  ;
  wire                xbar_mg3_ro_to_sg4_rsp_valid  ;
  wire                xbar_mg3_ro_to_sg4_rsp_err    ;
  wire                xbar_mg3_ro_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_ro_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg4_rsp_usr    ;
              wire                xbar_mg3_wo_to_sg4_cmd_valid  ;
  wire                xbar_mg3_wo_to_sg4_cmd_ready  ;
  wire                xbar_mg3_wo_to_sg4_cmd_sel    ;
  wire                xbar_mg3_wo_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg3_wo_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_wo_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_wo_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg4_cmd_size   ;
  wire                xbar_mg3_wo_to_sg4_cmd_lock   ;
  wire                xbar_mg3_wo_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_wo_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_wo_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_wo_to_sg4_cmd_modes  ;
  wire                xbar_mg3_wo_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_wo_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_wo_to_sg4_cmd_usr    ;
  wire                xbar_mg3_wo_to_sg4_rsp_ready  ;
  wire                xbar_mg3_wo_to_sg4_rsp_valid  ;
  wire                xbar_mg3_wo_to_sg4_rsp_err    ;
  wire                xbar_mg3_wo_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_wo_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg4_rsp_usr    ;
              wire                xbar_mg3_ro_to_sg5_cmd_valid  ;
  wire                xbar_mg3_ro_to_sg5_cmd_ready  ;
  wire                xbar_mg3_ro_to_sg5_cmd_sel    ;
  wire                xbar_mg3_ro_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg3_ro_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_ro_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_ro_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg5_cmd_size   ;
  wire                xbar_mg3_ro_to_sg5_cmd_lock   ;
  wire                xbar_mg3_ro_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_ro_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_ro_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_ro_to_sg5_cmd_modes  ;
  wire                xbar_mg3_ro_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_ro_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_ro_to_sg5_cmd_usr    ;
  wire                xbar_mg3_ro_to_sg5_rsp_ready  ;
  wire                xbar_mg3_ro_to_sg5_rsp_valid  ;
  wire                xbar_mg3_ro_to_sg5_rsp_err    ;
  wire                xbar_mg3_ro_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_ro_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg5_rsp_usr    ;
              wire                xbar_mg3_wo_to_sg5_cmd_valid  ;
  wire                xbar_mg3_wo_to_sg5_cmd_ready  ;
  wire                xbar_mg3_wo_to_sg5_cmd_sel    ;
  wire                xbar_mg3_wo_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg3_wo_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_wo_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_wo_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg5_cmd_size   ;
  wire                xbar_mg3_wo_to_sg5_cmd_lock   ;
  wire                xbar_mg3_wo_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_wo_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_wo_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_wo_to_sg5_cmd_modes  ;
  wire                xbar_mg3_wo_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_wo_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_wo_to_sg5_cmd_usr    ;
  wire                xbar_mg3_wo_to_sg5_rsp_ready  ;
  wire                xbar_mg3_wo_to_sg5_rsp_valid  ;
  wire                xbar_mg3_wo_to_sg5_rsp_err    ;
  wire                xbar_mg3_wo_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_wo_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg5_rsp_usr    ;
              wire                xbar_mg3_ro_to_sg6_cmd_valid  ;
  wire                xbar_mg3_ro_to_sg6_cmd_ready  ;
  wire                xbar_mg3_ro_to_sg6_cmd_sel    ;
  wire                xbar_mg3_ro_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg3_ro_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_ro_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_ro_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg6_cmd_size   ;
  wire                xbar_mg3_ro_to_sg6_cmd_lock   ;
  wire                xbar_mg3_ro_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_ro_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_ro_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_ro_to_sg6_cmd_modes  ;
  wire                xbar_mg3_ro_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_ro_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_ro_to_sg6_cmd_usr    ;
  wire                xbar_mg3_ro_to_sg6_rsp_ready  ;
  wire                xbar_mg3_ro_to_sg6_rsp_valid  ;
  wire                xbar_mg3_ro_to_sg6_rsp_err    ;
  wire                xbar_mg3_ro_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_ro_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_ro_to_sg6_rsp_usr    ;
              wire                xbar_mg3_wo_to_sg6_cmd_valid  ;
  wire                xbar_mg3_wo_to_sg6_cmd_ready  ;
  wire                xbar_mg3_wo_to_sg6_cmd_sel    ;
  wire                xbar_mg3_wo_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg3_wo_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg3_wo_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg3_wo_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg6_cmd_size   ;
  wire                xbar_mg3_wo_to_sg6_cmd_lock   ;
  wire                xbar_mg3_wo_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg3_wo_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg3_wo_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg3_wo_to_sg6_cmd_modes  ;
  wire                xbar_mg3_wo_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg3_wo_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg3_wo_to_sg6_cmd_usr    ;
  wire                xbar_mg3_wo_to_sg6_rsp_ready  ;
  wire                xbar_mg3_wo_to_sg6_rsp_valid  ;
  wire                xbar_mg3_wo_to_sg6_rsp_err    ;
  wire                xbar_mg3_wo_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg3_wo_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg3_wo_to_sg6_rsp_usr    ;
              wire                xbar_mg4_ro_to_sg0_cmd_valid  ;
  wire                xbar_mg4_ro_to_sg0_cmd_ready  ;
  wire                xbar_mg4_ro_to_sg0_cmd_sel    ;
  wire                xbar_mg4_ro_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg4_ro_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_ro_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_ro_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg0_cmd_size   ;
  wire                xbar_mg4_ro_to_sg0_cmd_lock   ;
  wire                xbar_mg4_ro_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_ro_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_ro_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_ro_to_sg0_cmd_modes  ;
  wire                xbar_mg4_ro_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_ro_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_ro_to_sg0_cmd_usr    ;
  wire                xbar_mg4_ro_to_sg0_rsp_ready  ;
  wire                xbar_mg4_ro_to_sg0_rsp_valid  ;
  wire                xbar_mg4_ro_to_sg0_rsp_err    ;
  wire                xbar_mg4_ro_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_ro_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg0_rsp_usr    ;
              wire                xbar_mg4_wo_to_sg0_cmd_valid  ;
  wire                xbar_mg4_wo_to_sg0_cmd_ready  ;
  wire                xbar_mg4_wo_to_sg0_cmd_sel    ;
  wire                xbar_mg4_wo_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg4_wo_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_wo_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_wo_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg0_cmd_size   ;
  wire                xbar_mg4_wo_to_sg0_cmd_lock   ;
  wire                xbar_mg4_wo_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_wo_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_wo_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_wo_to_sg0_cmd_modes  ;
  wire                xbar_mg4_wo_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_wo_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_wo_to_sg0_cmd_usr    ;
  wire                xbar_mg4_wo_to_sg0_rsp_ready  ;
  wire                xbar_mg4_wo_to_sg0_rsp_valid  ;
  wire                xbar_mg4_wo_to_sg0_rsp_err    ;
  wire                xbar_mg4_wo_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_wo_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg0_rsp_usr    ;
              wire                xbar_mg4_ro_to_sg1_cmd_valid  ;
  wire                xbar_mg4_ro_to_sg1_cmd_ready  ;
  wire                xbar_mg4_ro_to_sg1_cmd_sel    ;
  wire                xbar_mg4_ro_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg4_ro_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_ro_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_ro_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg1_cmd_size   ;
  wire                xbar_mg4_ro_to_sg1_cmd_lock   ;
  wire                xbar_mg4_ro_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_ro_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_ro_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_ro_to_sg1_cmd_modes  ;
  wire                xbar_mg4_ro_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_ro_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_ro_to_sg1_cmd_usr    ;
  wire                xbar_mg4_ro_to_sg1_rsp_ready  ;
  wire                xbar_mg4_ro_to_sg1_rsp_valid  ;
  wire                xbar_mg4_ro_to_sg1_rsp_err    ;
  wire                xbar_mg4_ro_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_ro_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg1_rsp_usr    ;
              wire                xbar_mg4_wo_to_sg1_cmd_valid  ;
  wire                xbar_mg4_wo_to_sg1_cmd_ready  ;
  wire                xbar_mg4_wo_to_sg1_cmd_sel    ;
  wire                xbar_mg4_wo_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg4_wo_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_wo_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_wo_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg1_cmd_size   ;
  wire                xbar_mg4_wo_to_sg1_cmd_lock   ;
  wire                xbar_mg4_wo_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_wo_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_wo_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_wo_to_sg1_cmd_modes  ;
  wire                xbar_mg4_wo_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_wo_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_wo_to_sg1_cmd_usr    ;
  wire                xbar_mg4_wo_to_sg1_rsp_ready  ;
  wire                xbar_mg4_wo_to_sg1_rsp_valid  ;
  wire                xbar_mg4_wo_to_sg1_rsp_err    ;
  wire                xbar_mg4_wo_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_wo_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg1_rsp_usr    ;
              wire                xbar_mg4_ro_to_sg2_cmd_valid  ;
  wire                xbar_mg4_ro_to_sg2_cmd_ready  ;
  wire                xbar_mg4_ro_to_sg2_cmd_sel    ;
  wire                xbar_mg4_ro_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg4_ro_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_ro_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_ro_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg2_cmd_size   ;
  wire                xbar_mg4_ro_to_sg2_cmd_lock   ;
  wire                xbar_mg4_ro_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_ro_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_ro_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_ro_to_sg2_cmd_modes  ;
  wire                xbar_mg4_ro_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_ro_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_ro_to_sg2_cmd_usr    ;
  wire                xbar_mg4_ro_to_sg2_rsp_ready  ;
  wire                xbar_mg4_ro_to_sg2_rsp_valid  ;
  wire                xbar_mg4_ro_to_sg2_rsp_err    ;
  wire                xbar_mg4_ro_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_ro_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg2_rsp_usr    ;
              wire                xbar_mg4_wo_to_sg2_cmd_valid  ;
  wire                xbar_mg4_wo_to_sg2_cmd_ready  ;
  wire                xbar_mg4_wo_to_sg2_cmd_sel    ;
  wire                xbar_mg4_wo_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg4_wo_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_wo_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_wo_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg2_cmd_size   ;
  wire                xbar_mg4_wo_to_sg2_cmd_lock   ;
  wire                xbar_mg4_wo_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_wo_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_wo_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_wo_to_sg2_cmd_modes  ;
  wire                xbar_mg4_wo_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_wo_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_wo_to_sg2_cmd_usr    ;
  wire                xbar_mg4_wo_to_sg2_rsp_ready  ;
  wire                xbar_mg4_wo_to_sg2_rsp_valid  ;
  wire                xbar_mg4_wo_to_sg2_rsp_err    ;
  wire                xbar_mg4_wo_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_wo_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg2_rsp_usr    ;
              wire                xbar_mg4_ro_to_sg3_cmd_valid  ;
  wire                xbar_mg4_ro_to_sg3_cmd_ready  ;
  wire                xbar_mg4_ro_to_sg3_cmd_sel    ;
  wire                xbar_mg4_ro_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg4_ro_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_ro_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_ro_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg3_cmd_size   ;
  wire                xbar_mg4_ro_to_sg3_cmd_lock   ;
  wire                xbar_mg4_ro_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_ro_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_ro_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_ro_to_sg3_cmd_modes  ;
  wire                xbar_mg4_ro_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_ro_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_ro_to_sg3_cmd_usr    ;
  wire                xbar_mg4_ro_to_sg3_rsp_ready  ;
  wire                xbar_mg4_ro_to_sg3_rsp_valid  ;
  wire                xbar_mg4_ro_to_sg3_rsp_err    ;
  wire                xbar_mg4_ro_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_ro_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg3_rsp_usr    ;
              wire                xbar_mg4_wo_to_sg3_cmd_valid  ;
  wire                xbar_mg4_wo_to_sg3_cmd_ready  ;
  wire                xbar_mg4_wo_to_sg3_cmd_sel    ;
  wire                xbar_mg4_wo_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg4_wo_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_wo_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_wo_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg3_cmd_size   ;
  wire                xbar_mg4_wo_to_sg3_cmd_lock   ;
  wire                xbar_mg4_wo_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_wo_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_wo_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_wo_to_sg3_cmd_modes  ;
  wire                xbar_mg4_wo_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_wo_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_wo_to_sg3_cmd_usr    ;
  wire                xbar_mg4_wo_to_sg3_rsp_ready  ;
  wire                xbar_mg4_wo_to_sg3_rsp_valid  ;
  wire                xbar_mg4_wo_to_sg3_rsp_err    ;
  wire                xbar_mg4_wo_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_wo_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg3_rsp_usr    ;
              wire                xbar_mg4_ro_to_sg4_cmd_valid  ;
  wire                xbar_mg4_ro_to_sg4_cmd_ready  ;
  wire                xbar_mg4_ro_to_sg4_cmd_sel    ;
  wire                xbar_mg4_ro_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg4_ro_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_ro_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_ro_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg4_cmd_size   ;
  wire                xbar_mg4_ro_to_sg4_cmd_lock   ;
  wire                xbar_mg4_ro_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_ro_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_ro_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_ro_to_sg4_cmd_modes  ;
  wire                xbar_mg4_ro_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_ro_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_ro_to_sg4_cmd_usr    ;
  wire                xbar_mg4_ro_to_sg4_rsp_ready  ;
  wire                xbar_mg4_ro_to_sg4_rsp_valid  ;
  wire                xbar_mg4_ro_to_sg4_rsp_err    ;
  wire                xbar_mg4_ro_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_ro_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg4_rsp_usr    ;
              wire                xbar_mg4_wo_to_sg4_cmd_valid  ;
  wire                xbar_mg4_wo_to_sg4_cmd_ready  ;
  wire                xbar_mg4_wo_to_sg4_cmd_sel    ;
  wire                xbar_mg4_wo_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg4_wo_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_wo_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_wo_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg4_cmd_size   ;
  wire                xbar_mg4_wo_to_sg4_cmd_lock   ;
  wire                xbar_mg4_wo_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_wo_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_wo_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_wo_to_sg4_cmd_modes  ;
  wire                xbar_mg4_wo_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_wo_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_wo_to_sg4_cmd_usr    ;
  wire                xbar_mg4_wo_to_sg4_rsp_ready  ;
  wire                xbar_mg4_wo_to_sg4_rsp_valid  ;
  wire                xbar_mg4_wo_to_sg4_rsp_err    ;
  wire                xbar_mg4_wo_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_wo_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg4_rsp_usr    ;
              wire                xbar_mg4_ro_to_sg5_cmd_valid  ;
  wire                xbar_mg4_ro_to_sg5_cmd_ready  ;
  wire                xbar_mg4_ro_to_sg5_cmd_sel    ;
  wire                xbar_mg4_ro_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg4_ro_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_ro_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_ro_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg5_cmd_size   ;
  wire                xbar_mg4_ro_to_sg5_cmd_lock   ;
  wire                xbar_mg4_ro_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_ro_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_ro_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_ro_to_sg5_cmd_modes  ;
  wire                xbar_mg4_ro_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_ro_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_ro_to_sg5_cmd_usr    ;
  wire                xbar_mg4_ro_to_sg5_rsp_ready  ;
  wire                xbar_mg4_ro_to_sg5_rsp_valid  ;
  wire                xbar_mg4_ro_to_sg5_rsp_err    ;
  wire                xbar_mg4_ro_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_ro_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg5_rsp_usr    ;
              wire                xbar_mg4_wo_to_sg5_cmd_valid  ;
  wire                xbar_mg4_wo_to_sg5_cmd_ready  ;
  wire                xbar_mg4_wo_to_sg5_cmd_sel    ;
  wire                xbar_mg4_wo_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg4_wo_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_wo_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_wo_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg5_cmd_size   ;
  wire                xbar_mg4_wo_to_sg5_cmd_lock   ;
  wire                xbar_mg4_wo_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_wo_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_wo_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_wo_to_sg5_cmd_modes  ;
  wire                xbar_mg4_wo_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_wo_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_wo_to_sg5_cmd_usr    ;
  wire                xbar_mg4_wo_to_sg5_rsp_ready  ;
  wire                xbar_mg4_wo_to_sg5_rsp_valid  ;
  wire                xbar_mg4_wo_to_sg5_rsp_err    ;
  wire                xbar_mg4_wo_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_wo_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg5_rsp_usr    ;
              wire                xbar_mg4_ro_to_sg6_cmd_valid  ;
  wire                xbar_mg4_ro_to_sg6_cmd_ready  ;
  wire                xbar_mg4_ro_to_sg6_cmd_sel    ;
  wire                xbar_mg4_ro_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg4_ro_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_ro_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_ro_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg6_cmd_size   ;
  wire                xbar_mg4_ro_to_sg6_cmd_lock   ;
  wire                xbar_mg4_ro_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_ro_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_ro_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_ro_to_sg6_cmd_modes  ;
  wire                xbar_mg4_ro_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_ro_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_ro_to_sg6_cmd_usr    ;
  wire                xbar_mg4_ro_to_sg6_rsp_ready  ;
  wire                xbar_mg4_ro_to_sg6_rsp_valid  ;
  wire                xbar_mg4_ro_to_sg6_rsp_err    ;
  wire                xbar_mg4_ro_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_ro_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_ro_to_sg6_rsp_usr    ;
              wire                xbar_mg4_wo_to_sg6_cmd_valid  ;
  wire                xbar_mg4_wo_to_sg6_cmd_ready  ;
  wire                xbar_mg4_wo_to_sg6_cmd_sel    ;
  wire                xbar_mg4_wo_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg4_wo_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg4_wo_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg4_wo_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg6_cmd_size   ;
  wire                xbar_mg4_wo_to_sg6_cmd_lock   ;
  wire                xbar_mg4_wo_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg4_wo_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg4_wo_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg4_wo_to_sg6_cmd_modes  ;
  wire                xbar_mg4_wo_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg4_wo_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg4_wo_to_sg6_cmd_usr    ;
  wire                xbar_mg4_wo_to_sg6_rsp_ready  ;
  wire                xbar_mg4_wo_to_sg6_rsp_valid  ;
  wire                xbar_mg4_wo_to_sg6_rsp_err    ;
  wire                xbar_mg4_wo_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg4_wo_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg4_wo_to_sg6_rsp_usr    ;
              wire                xbar_mg5_ro_to_sg0_cmd_valid  ;
  wire                xbar_mg5_ro_to_sg0_cmd_ready  ;
  wire                xbar_mg5_ro_to_sg0_cmd_sel    ;
  wire                xbar_mg5_ro_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg5_ro_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_ro_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_ro_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg0_cmd_size   ;
  wire                xbar_mg5_ro_to_sg0_cmd_lock   ;
  wire                xbar_mg5_ro_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_ro_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_ro_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_ro_to_sg0_cmd_modes  ;
  wire                xbar_mg5_ro_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_ro_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_ro_to_sg0_cmd_usr    ;
  wire                xbar_mg5_ro_to_sg0_rsp_ready  ;
  wire                xbar_mg5_ro_to_sg0_rsp_valid  ;
  wire                xbar_mg5_ro_to_sg0_rsp_err    ;
  wire                xbar_mg5_ro_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_ro_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg0_rsp_usr    ;
              wire                xbar_mg5_wo_to_sg0_cmd_valid  ;
  wire                xbar_mg5_wo_to_sg0_cmd_ready  ;
  wire                xbar_mg5_wo_to_sg0_cmd_sel    ;
  wire                xbar_mg5_wo_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg5_wo_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_wo_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_wo_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg0_cmd_size   ;
  wire                xbar_mg5_wo_to_sg0_cmd_lock   ;
  wire                xbar_mg5_wo_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_wo_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_wo_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_wo_to_sg0_cmd_modes  ;
  wire                xbar_mg5_wo_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_wo_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_wo_to_sg0_cmd_usr    ;
  wire                xbar_mg5_wo_to_sg0_rsp_ready  ;
  wire                xbar_mg5_wo_to_sg0_rsp_valid  ;
  wire                xbar_mg5_wo_to_sg0_rsp_err    ;
  wire                xbar_mg5_wo_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_wo_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg0_rsp_usr    ;
              wire                xbar_mg5_ro_to_sg1_cmd_valid  ;
  wire                xbar_mg5_ro_to_sg1_cmd_ready  ;
  wire                xbar_mg5_ro_to_sg1_cmd_sel    ;
  wire                xbar_mg5_ro_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg5_ro_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_ro_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_ro_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg1_cmd_size   ;
  wire                xbar_mg5_ro_to_sg1_cmd_lock   ;
  wire                xbar_mg5_ro_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_ro_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_ro_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_ro_to_sg1_cmd_modes  ;
  wire                xbar_mg5_ro_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_ro_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_ro_to_sg1_cmd_usr    ;
  wire                xbar_mg5_ro_to_sg1_rsp_ready  ;
  wire                xbar_mg5_ro_to_sg1_rsp_valid  ;
  wire                xbar_mg5_ro_to_sg1_rsp_err    ;
  wire                xbar_mg5_ro_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_ro_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg1_rsp_usr    ;
              wire                xbar_mg5_wo_to_sg1_cmd_valid  ;
  wire                xbar_mg5_wo_to_sg1_cmd_ready  ;
  wire                xbar_mg5_wo_to_sg1_cmd_sel    ;
  wire                xbar_mg5_wo_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg5_wo_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_wo_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_wo_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg1_cmd_size   ;
  wire                xbar_mg5_wo_to_sg1_cmd_lock   ;
  wire                xbar_mg5_wo_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_wo_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_wo_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_wo_to_sg1_cmd_modes  ;
  wire                xbar_mg5_wo_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_wo_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_wo_to_sg1_cmd_usr    ;
  wire                xbar_mg5_wo_to_sg1_rsp_ready  ;
  wire                xbar_mg5_wo_to_sg1_rsp_valid  ;
  wire                xbar_mg5_wo_to_sg1_rsp_err    ;
  wire                xbar_mg5_wo_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_wo_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg1_rsp_usr    ;
              wire                xbar_mg5_ro_to_sg2_cmd_valid  ;
  wire                xbar_mg5_ro_to_sg2_cmd_ready  ;
  wire                xbar_mg5_ro_to_sg2_cmd_sel    ;
  wire                xbar_mg5_ro_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg5_ro_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_ro_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_ro_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg2_cmd_size   ;
  wire                xbar_mg5_ro_to_sg2_cmd_lock   ;
  wire                xbar_mg5_ro_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_ro_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_ro_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_ro_to_sg2_cmd_modes  ;
  wire                xbar_mg5_ro_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_ro_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_ro_to_sg2_cmd_usr    ;
  wire                xbar_mg5_ro_to_sg2_rsp_ready  ;
  wire                xbar_mg5_ro_to_sg2_rsp_valid  ;
  wire                xbar_mg5_ro_to_sg2_rsp_err    ;
  wire                xbar_mg5_ro_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_ro_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg2_rsp_usr    ;
              wire                xbar_mg5_wo_to_sg2_cmd_valid  ;
  wire                xbar_mg5_wo_to_sg2_cmd_ready  ;
  wire                xbar_mg5_wo_to_sg2_cmd_sel    ;
  wire                xbar_mg5_wo_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg5_wo_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_wo_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_wo_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg2_cmd_size   ;
  wire                xbar_mg5_wo_to_sg2_cmd_lock   ;
  wire                xbar_mg5_wo_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_wo_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_wo_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_wo_to_sg2_cmd_modes  ;
  wire                xbar_mg5_wo_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_wo_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_wo_to_sg2_cmd_usr    ;
  wire                xbar_mg5_wo_to_sg2_rsp_ready  ;
  wire                xbar_mg5_wo_to_sg2_rsp_valid  ;
  wire                xbar_mg5_wo_to_sg2_rsp_err    ;
  wire                xbar_mg5_wo_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_wo_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg2_rsp_usr    ;
              wire                xbar_mg5_ro_to_sg3_cmd_valid  ;
  wire                xbar_mg5_ro_to_sg3_cmd_ready  ;
  wire                xbar_mg5_ro_to_sg3_cmd_sel    ;
  wire                xbar_mg5_ro_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg5_ro_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_ro_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_ro_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg3_cmd_size   ;
  wire                xbar_mg5_ro_to_sg3_cmd_lock   ;
  wire                xbar_mg5_ro_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_ro_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_ro_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_ro_to_sg3_cmd_modes  ;
  wire                xbar_mg5_ro_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_ro_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_ro_to_sg3_cmd_usr    ;
  wire                xbar_mg5_ro_to_sg3_rsp_ready  ;
  wire                xbar_mg5_ro_to_sg3_rsp_valid  ;
  wire                xbar_mg5_ro_to_sg3_rsp_err    ;
  wire                xbar_mg5_ro_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_ro_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg3_rsp_usr    ;
              wire                xbar_mg5_wo_to_sg3_cmd_valid  ;
  wire                xbar_mg5_wo_to_sg3_cmd_ready  ;
  wire                xbar_mg5_wo_to_sg3_cmd_sel    ;
  wire                xbar_mg5_wo_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg5_wo_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_wo_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_wo_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg3_cmd_size   ;
  wire                xbar_mg5_wo_to_sg3_cmd_lock   ;
  wire                xbar_mg5_wo_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_wo_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_wo_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_wo_to_sg3_cmd_modes  ;
  wire                xbar_mg5_wo_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_wo_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_wo_to_sg3_cmd_usr    ;
  wire                xbar_mg5_wo_to_sg3_rsp_ready  ;
  wire                xbar_mg5_wo_to_sg3_rsp_valid  ;
  wire                xbar_mg5_wo_to_sg3_rsp_err    ;
  wire                xbar_mg5_wo_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_wo_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg3_rsp_usr    ;
              wire                xbar_mg5_ro_to_sg4_cmd_valid  ;
  wire                xbar_mg5_ro_to_sg4_cmd_ready  ;
  wire                xbar_mg5_ro_to_sg4_cmd_sel    ;
  wire                xbar_mg5_ro_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg5_ro_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_ro_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_ro_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg4_cmd_size   ;
  wire                xbar_mg5_ro_to_sg4_cmd_lock   ;
  wire                xbar_mg5_ro_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_ro_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_ro_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_ro_to_sg4_cmd_modes  ;
  wire                xbar_mg5_ro_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_ro_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_ro_to_sg4_cmd_usr    ;
  wire                xbar_mg5_ro_to_sg4_rsp_ready  ;
  wire                xbar_mg5_ro_to_sg4_rsp_valid  ;
  wire                xbar_mg5_ro_to_sg4_rsp_err    ;
  wire                xbar_mg5_ro_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_ro_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg4_rsp_usr    ;
              wire                xbar_mg5_wo_to_sg4_cmd_valid  ;
  wire                xbar_mg5_wo_to_sg4_cmd_ready  ;
  wire                xbar_mg5_wo_to_sg4_cmd_sel    ;
  wire                xbar_mg5_wo_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg5_wo_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_wo_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_wo_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg4_cmd_size   ;
  wire                xbar_mg5_wo_to_sg4_cmd_lock   ;
  wire                xbar_mg5_wo_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_wo_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_wo_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_wo_to_sg4_cmd_modes  ;
  wire                xbar_mg5_wo_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_wo_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_wo_to_sg4_cmd_usr    ;
  wire                xbar_mg5_wo_to_sg4_rsp_ready  ;
  wire                xbar_mg5_wo_to_sg4_rsp_valid  ;
  wire                xbar_mg5_wo_to_sg4_rsp_err    ;
  wire                xbar_mg5_wo_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_wo_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg4_rsp_usr    ;
              wire                xbar_mg5_ro_to_sg5_cmd_valid  ;
  wire                xbar_mg5_ro_to_sg5_cmd_ready  ;
  wire                xbar_mg5_ro_to_sg5_cmd_sel    ;
  wire                xbar_mg5_ro_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg5_ro_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_ro_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_ro_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg5_cmd_size   ;
  wire                xbar_mg5_ro_to_sg5_cmd_lock   ;
  wire                xbar_mg5_ro_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_ro_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_ro_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_ro_to_sg5_cmd_modes  ;
  wire                xbar_mg5_ro_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_ro_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_ro_to_sg5_cmd_usr    ;
  wire                xbar_mg5_ro_to_sg5_rsp_ready  ;
  wire                xbar_mg5_ro_to_sg5_rsp_valid  ;
  wire                xbar_mg5_ro_to_sg5_rsp_err    ;
  wire                xbar_mg5_ro_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_ro_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg5_rsp_usr    ;
              wire                xbar_mg5_wo_to_sg5_cmd_valid  ;
  wire                xbar_mg5_wo_to_sg5_cmd_ready  ;
  wire                xbar_mg5_wo_to_sg5_cmd_sel    ;
  wire                xbar_mg5_wo_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg5_wo_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_wo_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_wo_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg5_cmd_size   ;
  wire                xbar_mg5_wo_to_sg5_cmd_lock   ;
  wire                xbar_mg5_wo_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_wo_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_wo_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_wo_to_sg5_cmd_modes  ;
  wire                xbar_mg5_wo_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_wo_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_wo_to_sg5_cmd_usr    ;
  wire                xbar_mg5_wo_to_sg5_rsp_ready  ;
  wire                xbar_mg5_wo_to_sg5_rsp_valid  ;
  wire                xbar_mg5_wo_to_sg5_rsp_err    ;
  wire                xbar_mg5_wo_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_wo_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg5_rsp_usr    ;
              wire                xbar_mg5_ro_to_sg6_cmd_valid  ;
  wire                xbar_mg5_ro_to_sg6_cmd_ready  ;
  wire                xbar_mg5_ro_to_sg6_cmd_sel    ;
  wire                xbar_mg5_ro_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg5_ro_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_ro_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_ro_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg6_cmd_size   ;
  wire                xbar_mg5_ro_to_sg6_cmd_lock   ;
  wire                xbar_mg5_ro_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_ro_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_ro_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_ro_to_sg6_cmd_modes  ;
  wire                xbar_mg5_ro_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_ro_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_ro_to_sg6_cmd_usr    ;
  wire                xbar_mg5_ro_to_sg6_rsp_ready  ;
  wire                xbar_mg5_ro_to_sg6_rsp_valid  ;
  wire                xbar_mg5_ro_to_sg6_rsp_err    ;
  wire                xbar_mg5_ro_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_ro_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_ro_to_sg6_rsp_usr    ;
              wire                xbar_mg5_wo_to_sg6_cmd_valid  ;
  wire                xbar_mg5_wo_to_sg6_cmd_ready  ;
  wire                xbar_mg5_wo_to_sg6_cmd_sel    ;
  wire                xbar_mg5_wo_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg5_wo_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg5_wo_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg5_wo_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg6_cmd_size   ;
  wire                xbar_mg5_wo_to_sg6_cmd_lock   ;
  wire                xbar_mg5_wo_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg5_wo_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg5_wo_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg5_wo_to_sg6_cmd_modes  ;
  wire                xbar_mg5_wo_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg5_wo_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg5_wo_to_sg6_cmd_usr    ;
  wire                xbar_mg5_wo_to_sg6_rsp_ready  ;
  wire                xbar_mg5_wo_to_sg6_rsp_valid  ;
  wire                xbar_mg5_wo_to_sg6_rsp_err    ;
  wire                xbar_mg5_wo_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg5_wo_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg5_wo_to_sg6_rsp_usr    ;
              wire                xbar_mg6_ro_to_sg0_cmd_valid  ;
  wire                xbar_mg6_ro_to_sg0_cmd_ready  ;
  wire                xbar_mg6_ro_to_sg0_cmd_sel    ;
  wire                xbar_mg6_ro_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg6_ro_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_ro_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_ro_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg0_cmd_size   ;
  wire                xbar_mg6_ro_to_sg0_cmd_lock   ;
  wire                xbar_mg6_ro_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_ro_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_ro_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_ro_to_sg0_cmd_modes  ;
  wire                xbar_mg6_ro_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_ro_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_ro_to_sg0_cmd_usr    ;
  wire                xbar_mg6_ro_to_sg0_rsp_ready  ;
  wire                xbar_mg6_ro_to_sg0_rsp_valid  ;
  wire                xbar_mg6_ro_to_sg0_rsp_err    ;
  wire                xbar_mg6_ro_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_ro_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg0_rsp_usr    ;
              wire                xbar_mg6_wo_to_sg0_cmd_valid  ;
  wire                xbar_mg6_wo_to_sg0_cmd_ready  ;
  wire                xbar_mg6_wo_to_sg0_cmd_sel    ;
  wire                xbar_mg6_wo_to_sg0_cmd_read   ;
  wire    [  31:   0] xbar_mg6_wo_to_sg0_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_wo_to_sg0_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_wo_to_sg0_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg0_cmd_size   ;
  wire                xbar_mg6_wo_to_sg0_cmd_lock   ;
  wire                xbar_mg6_wo_to_sg0_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_wo_to_sg0_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_wo_to_sg0_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_wo_to_sg0_cmd_modes  ;
  wire                xbar_mg6_wo_to_sg0_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg0_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_wo_to_sg0_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_wo_to_sg0_cmd_usr    ;
  wire                xbar_mg6_wo_to_sg0_rsp_ready  ;
  wire                xbar_mg6_wo_to_sg0_rsp_valid  ;
  wire                xbar_mg6_wo_to_sg0_rsp_err    ;
  wire                xbar_mg6_wo_to_sg0_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_wo_to_sg0_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg0_rsp_usr    ;
              wire                xbar_mg6_ro_to_sg1_cmd_valid  ;
  wire                xbar_mg6_ro_to_sg1_cmd_ready  ;
  wire                xbar_mg6_ro_to_sg1_cmd_sel    ;
  wire                xbar_mg6_ro_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg6_ro_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_ro_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_ro_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg1_cmd_size   ;
  wire                xbar_mg6_ro_to_sg1_cmd_lock   ;
  wire                xbar_mg6_ro_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_ro_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_ro_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_ro_to_sg1_cmd_modes  ;
  wire                xbar_mg6_ro_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_ro_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_ro_to_sg1_cmd_usr    ;
  wire                xbar_mg6_ro_to_sg1_rsp_ready  ;
  wire                xbar_mg6_ro_to_sg1_rsp_valid  ;
  wire                xbar_mg6_ro_to_sg1_rsp_err    ;
  wire                xbar_mg6_ro_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_ro_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg1_rsp_usr    ;
              wire                xbar_mg6_wo_to_sg1_cmd_valid  ;
  wire                xbar_mg6_wo_to_sg1_cmd_ready  ;
  wire                xbar_mg6_wo_to_sg1_cmd_sel    ;
  wire                xbar_mg6_wo_to_sg1_cmd_read   ;
  wire    [  31:   0] xbar_mg6_wo_to_sg1_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_wo_to_sg1_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_wo_to_sg1_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg1_cmd_size   ;
  wire                xbar_mg6_wo_to_sg1_cmd_lock   ;
  wire                xbar_mg6_wo_to_sg1_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_wo_to_sg1_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_wo_to_sg1_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_wo_to_sg1_cmd_modes  ;
  wire                xbar_mg6_wo_to_sg1_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg1_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_wo_to_sg1_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_wo_to_sg1_cmd_usr    ;
  wire                xbar_mg6_wo_to_sg1_rsp_ready  ;
  wire                xbar_mg6_wo_to_sg1_rsp_valid  ;
  wire                xbar_mg6_wo_to_sg1_rsp_err    ;
  wire                xbar_mg6_wo_to_sg1_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_wo_to_sg1_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg1_rsp_usr    ;
              wire                xbar_mg6_ro_to_sg2_cmd_valid  ;
  wire                xbar_mg6_ro_to_sg2_cmd_ready  ;
  wire                xbar_mg6_ro_to_sg2_cmd_sel    ;
  wire                xbar_mg6_ro_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg6_ro_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_ro_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_ro_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg2_cmd_size   ;
  wire                xbar_mg6_ro_to_sg2_cmd_lock   ;
  wire                xbar_mg6_ro_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_ro_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_ro_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_ro_to_sg2_cmd_modes  ;
  wire                xbar_mg6_ro_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_ro_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_ro_to_sg2_cmd_usr    ;
  wire                xbar_mg6_ro_to_sg2_rsp_ready  ;
  wire                xbar_mg6_ro_to_sg2_rsp_valid  ;
  wire                xbar_mg6_ro_to_sg2_rsp_err    ;
  wire                xbar_mg6_ro_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_ro_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg2_rsp_usr    ;
              wire                xbar_mg6_wo_to_sg2_cmd_valid  ;
  wire                xbar_mg6_wo_to_sg2_cmd_ready  ;
  wire                xbar_mg6_wo_to_sg2_cmd_sel    ;
  wire                xbar_mg6_wo_to_sg2_cmd_read   ;
  wire    [  31:   0] xbar_mg6_wo_to_sg2_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_wo_to_sg2_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_wo_to_sg2_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg2_cmd_size   ;
  wire                xbar_mg6_wo_to_sg2_cmd_lock   ;
  wire                xbar_mg6_wo_to_sg2_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_wo_to_sg2_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_wo_to_sg2_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_wo_to_sg2_cmd_modes  ;
  wire                xbar_mg6_wo_to_sg2_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg2_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_wo_to_sg2_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_wo_to_sg2_cmd_usr    ;
  wire                xbar_mg6_wo_to_sg2_rsp_ready  ;
  wire                xbar_mg6_wo_to_sg2_rsp_valid  ;
  wire                xbar_mg6_wo_to_sg2_rsp_err    ;
  wire                xbar_mg6_wo_to_sg2_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_wo_to_sg2_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg2_rsp_usr    ;
              wire                xbar_mg6_ro_to_sg3_cmd_valid  ;
  wire                xbar_mg6_ro_to_sg3_cmd_ready  ;
  wire                xbar_mg6_ro_to_sg3_cmd_sel    ;
  wire                xbar_mg6_ro_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg6_ro_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_ro_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_ro_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg3_cmd_size   ;
  wire                xbar_mg6_ro_to_sg3_cmd_lock   ;
  wire                xbar_mg6_ro_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_ro_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_ro_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_ro_to_sg3_cmd_modes  ;
  wire                xbar_mg6_ro_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_ro_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_ro_to_sg3_cmd_usr    ;
  wire                xbar_mg6_ro_to_sg3_rsp_ready  ;
  wire                xbar_mg6_ro_to_sg3_rsp_valid  ;
  wire                xbar_mg6_ro_to_sg3_rsp_err    ;
  wire                xbar_mg6_ro_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_ro_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg3_rsp_usr    ;
              wire                xbar_mg6_wo_to_sg3_cmd_valid  ;
  wire                xbar_mg6_wo_to_sg3_cmd_ready  ;
  wire                xbar_mg6_wo_to_sg3_cmd_sel    ;
  wire                xbar_mg6_wo_to_sg3_cmd_read   ;
  wire    [  31:   0] xbar_mg6_wo_to_sg3_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_wo_to_sg3_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_wo_to_sg3_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg3_cmd_size   ;
  wire                xbar_mg6_wo_to_sg3_cmd_lock   ;
  wire                xbar_mg6_wo_to_sg3_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_wo_to_sg3_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_wo_to_sg3_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_wo_to_sg3_cmd_modes  ;
  wire                xbar_mg6_wo_to_sg3_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg3_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_wo_to_sg3_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_wo_to_sg3_cmd_usr    ;
  wire                xbar_mg6_wo_to_sg3_rsp_ready  ;
  wire                xbar_mg6_wo_to_sg3_rsp_valid  ;
  wire                xbar_mg6_wo_to_sg3_rsp_err    ;
  wire                xbar_mg6_wo_to_sg3_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_wo_to_sg3_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg3_rsp_usr    ;
              wire                xbar_mg6_ro_to_sg4_cmd_valid  ;
  wire                xbar_mg6_ro_to_sg4_cmd_ready  ;
  wire                xbar_mg6_ro_to_sg4_cmd_sel    ;
  wire                xbar_mg6_ro_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg6_ro_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_ro_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_ro_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg4_cmd_size   ;
  wire                xbar_mg6_ro_to_sg4_cmd_lock   ;
  wire                xbar_mg6_ro_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_ro_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_ro_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_ro_to_sg4_cmd_modes  ;
  wire                xbar_mg6_ro_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_ro_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_ro_to_sg4_cmd_usr    ;
  wire                xbar_mg6_ro_to_sg4_rsp_ready  ;
  wire                xbar_mg6_ro_to_sg4_rsp_valid  ;
  wire                xbar_mg6_ro_to_sg4_rsp_err    ;
  wire                xbar_mg6_ro_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_ro_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg4_rsp_usr    ;
              wire                xbar_mg6_wo_to_sg4_cmd_valid  ;
  wire                xbar_mg6_wo_to_sg4_cmd_ready  ;
  wire                xbar_mg6_wo_to_sg4_cmd_sel    ;
  wire                xbar_mg6_wo_to_sg4_cmd_read   ;
  wire    [  31:   0] xbar_mg6_wo_to_sg4_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_wo_to_sg4_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_wo_to_sg4_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg4_cmd_size   ;
  wire                xbar_mg6_wo_to_sg4_cmd_lock   ;
  wire                xbar_mg6_wo_to_sg4_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_wo_to_sg4_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_wo_to_sg4_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_wo_to_sg4_cmd_modes  ;
  wire                xbar_mg6_wo_to_sg4_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg4_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_wo_to_sg4_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_wo_to_sg4_cmd_usr    ;
  wire                xbar_mg6_wo_to_sg4_rsp_ready  ;
  wire                xbar_mg6_wo_to_sg4_rsp_valid  ;
  wire                xbar_mg6_wo_to_sg4_rsp_err    ;
  wire                xbar_mg6_wo_to_sg4_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_wo_to_sg4_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg4_rsp_usr    ;
              wire                xbar_mg6_ro_to_sg5_cmd_valid  ;
  wire                xbar_mg6_ro_to_sg5_cmd_ready  ;
  wire                xbar_mg6_ro_to_sg5_cmd_sel    ;
  wire                xbar_mg6_ro_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg6_ro_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_ro_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_ro_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg5_cmd_size   ;
  wire                xbar_mg6_ro_to_sg5_cmd_lock   ;
  wire                xbar_mg6_ro_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_ro_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_ro_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_ro_to_sg5_cmd_modes  ;
  wire                xbar_mg6_ro_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_ro_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_ro_to_sg5_cmd_usr    ;
  wire                xbar_mg6_ro_to_sg5_rsp_ready  ;
  wire                xbar_mg6_ro_to_sg5_rsp_valid  ;
  wire                xbar_mg6_ro_to_sg5_rsp_err    ;
  wire                xbar_mg6_ro_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_ro_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg5_rsp_usr    ;
              wire                xbar_mg6_wo_to_sg5_cmd_valid  ;
  wire                xbar_mg6_wo_to_sg5_cmd_ready  ;
  wire                xbar_mg6_wo_to_sg5_cmd_sel    ;
  wire                xbar_mg6_wo_to_sg5_cmd_read   ;
  wire    [  31:   0] xbar_mg6_wo_to_sg5_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_wo_to_sg5_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_wo_to_sg5_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg5_cmd_size   ;
  wire                xbar_mg6_wo_to_sg5_cmd_lock   ;
  wire                xbar_mg6_wo_to_sg5_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_wo_to_sg5_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_wo_to_sg5_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_wo_to_sg5_cmd_modes  ;
  wire                xbar_mg6_wo_to_sg5_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg5_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_wo_to_sg5_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_wo_to_sg5_cmd_usr    ;
  wire                xbar_mg6_wo_to_sg5_rsp_ready  ;
  wire                xbar_mg6_wo_to_sg5_rsp_valid  ;
  wire                xbar_mg6_wo_to_sg5_rsp_err    ;
  wire                xbar_mg6_wo_to_sg5_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_wo_to_sg5_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg5_rsp_usr    ;
              wire                xbar_mg6_ro_to_sg6_cmd_valid  ;
  wire                xbar_mg6_ro_to_sg6_cmd_ready  ;
  wire                xbar_mg6_ro_to_sg6_cmd_sel    ;
  wire                xbar_mg6_ro_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg6_ro_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_ro_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_ro_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg6_cmd_size   ;
  wire                xbar_mg6_ro_to_sg6_cmd_lock   ;
  wire                xbar_mg6_ro_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_ro_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_ro_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_ro_to_sg6_cmd_modes  ;
  wire                xbar_mg6_ro_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_ro_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_ro_to_sg6_cmd_usr    ;
  wire                xbar_mg6_ro_to_sg6_rsp_ready  ;
  wire                xbar_mg6_ro_to_sg6_rsp_valid  ;
  wire                xbar_mg6_ro_to_sg6_rsp_err    ;
  wire                xbar_mg6_ro_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_ro_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_ro_to_sg6_rsp_usr    ;
              wire                xbar_mg6_wo_to_sg6_cmd_valid  ;
  wire                xbar_mg6_wo_to_sg6_cmd_ready  ;
  wire                xbar_mg6_wo_to_sg6_cmd_sel    ;
  wire                xbar_mg6_wo_to_sg6_cmd_read   ;
  wire    [  31:   0] xbar_mg6_wo_to_sg6_cmd_addr   ;
  wire    [  63:   0] xbar_mg6_wo_to_sg6_cmd_wdata  ;
  wire    [   7:   0] xbar_mg6_wo_to_sg6_cmd_wmask  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg6_cmd_size   ;
  wire                xbar_mg6_wo_to_sg6_cmd_lock   ;
  wire                xbar_mg6_wo_to_sg6_cmd_excl   ;
  wire    [   7:   0] xbar_mg6_wo_to_sg6_cmd_xlen   ;
  wire    [   1:   0] xbar_mg6_wo_to_sg6_cmd_xburst ;
  wire    [   1:   0] xbar_mg6_wo_to_sg6_cmd_modes  ;
  wire                xbar_mg6_wo_to_sg6_cmd_dmode  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg6_cmd_attri  ;
  wire    [   1:   0] xbar_mg6_wo_to_sg6_cmd_beat   ;
  wire    [   2:   0] xbar_mg6_wo_to_sg6_cmd_usr    ;
  wire                xbar_mg6_wo_to_sg6_rsp_ready  ;
  wire                xbar_mg6_wo_to_sg6_rsp_valid  ;
  wire                xbar_mg6_wo_to_sg6_rsp_err    ;
  wire                xbar_mg6_wo_to_sg6_rsp_excl_ok ;
  wire    [  63:   0] xbar_mg6_wo_to_sg6_rsp_rdata  ;
  wire    [   2:   0] xbar_mg6_wo_to_sg6_rsp_usr    ;
      wire                mst_grp_3_ro_icb_cmd_valid    ;
  wire                mst_grp_3_ro_icb_cmd_ready    ;
  wire                mst_grp_3_ro_icb_cmd_sel      ;
  wire                mst_grp_3_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_3_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_3_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_3_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_3_ro_icb_cmd_size     ;
  wire                mst_grp_3_ro_icb_cmd_lock     ;
  wire                mst_grp_3_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_3_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_3_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_3_ro_icb_cmd_modes    ;
  wire                mst_grp_3_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_3_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_3_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_3_ro_icb_cmd_usr      ;
  wire                mst_grp_3_ro_icb_rsp_ready    ;
  wire                mst_grp_3_ro_icb_rsp_valid    ;
  wire                mst_grp_3_ro_icb_rsp_err      ;
  wire                mst_grp_3_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_3_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_3_ro_icb_rsp_usr      ;
      wire                mst_grp_3_wo_icb_cmd_valid    ;
  wire                mst_grp_3_wo_icb_cmd_ready    ;
  wire                mst_grp_3_wo_icb_cmd_sel      ;
  wire                mst_grp_3_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_3_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_3_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_3_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_3_wo_icb_cmd_size     ;
  wire                mst_grp_3_wo_icb_cmd_lock     ;
  wire                mst_grp_3_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_3_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_3_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_3_wo_icb_cmd_modes    ;
  wire                mst_grp_3_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_3_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_3_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_3_wo_icb_cmd_usr      ;
  wire                mst_grp_3_wo_icb_rsp_ready    ;
  wire                mst_grp_3_wo_icb_rsp_valid    ;
  wire                mst_grp_3_wo_icb_rsp_err      ;
  wire                mst_grp_3_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_3_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_3_wo_icb_rsp_usr      ;
  e603_subsys_gnrl_ficb_rw_splt # (
      .ALLOW_DIFF   (0),
      .AW           (32),
      .DW           (64),
      .OUTS_FIFO_DP (64),
      .CMD_UW       (3),
      .RSP_UW       (3) 
   ) u_xbar_mg3_rw_splt(
      .icb_cmd_valid                  (mst_grp_3_icb_cmd_valid                  ),
  .icb_cmd_ready                  (mst_grp_3_icb_cmd_ready                  ),
  .icb_cmd_sel                    (mst_grp_3_icb_cmd_sel                    ),
  .icb_cmd_read                   (mst_grp_3_icb_cmd_read                   ),
  .icb_cmd_addr                   (mst_grp_3_icb_cmd_addr        [  31:   0]),
  .icb_cmd_wdata                  (mst_grp_3_icb_cmd_wdata       [  63:   0]),
  .icb_cmd_wmask                  (mst_grp_3_icb_cmd_wmask       [   7:   0]),
  .icb_cmd_size                   (mst_grp_3_icb_cmd_size        [   2:   0]),
  .icb_cmd_lock                   (mst_grp_3_icb_cmd_lock                   ),
  .icb_cmd_excl                   (mst_grp_3_icb_cmd_excl                   ),
  .icb_cmd_xlen                   (mst_grp_3_icb_cmd_xlen        [   7:   0]),
  .icb_cmd_xburst                 (mst_grp_3_icb_cmd_xburst      [   1:   0]),
  .icb_cmd_modes                  (mst_grp_3_icb_cmd_modes       [   1:   0]),
  .icb_cmd_dmode                  (mst_grp_3_icb_cmd_dmode                  ),
  .icb_cmd_attri                  (mst_grp_3_icb_cmd_attri       [   2:   0]),
  .icb_cmd_beat                   (mst_grp_3_icb_cmd_beat        [   1:   0]),
  .icb_cmd_usr                    (mst_grp_3_icb_cmd_usr         [   2:   0]),
  .icb_rsp_ready                  (mst_grp_3_icb_rsp_ready                  ),
  .icb_rsp_valid                  (mst_grp_3_icb_rsp_valid                  ),
  .icb_rsp_err                    (mst_grp_3_icb_rsp_err                    ),
  .icb_rsp_excl_ok                (mst_grp_3_icb_rsp_excl_ok                ),
  .icb_rsp_rdata                  (mst_grp_3_icb_rsp_rdata       [  63:   0]),
  .icb_rsp_usr                    (mst_grp_3_icb_rsp_usr         [   2:   0]),
      .r_icb_cmd_valid                (mst_grp_3_ro_icb_cmd_valid               ),
  .r_icb_cmd_ready                (mst_grp_3_ro_icb_cmd_ready               ),
  .r_icb_cmd_sel                  (mst_grp_3_ro_icb_cmd_sel                 ),
  .r_icb_cmd_read                 (mst_grp_3_ro_icb_cmd_read                ),
  .r_icb_cmd_addr                 (mst_grp_3_ro_icb_cmd_addr     [  31:   0]),
  .r_icb_cmd_wdata                (mst_grp_3_ro_icb_cmd_wdata    [  63:   0]),
  .r_icb_cmd_wmask                (mst_grp_3_ro_icb_cmd_wmask    [   7:   0]),
  .r_icb_cmd_size                 (mst_grp_3_ro_icb_cmd_size     [   2:   0]),
  .r_icb_cmd_lock                 (mst_grp_3_ro_icb_cmd_lock                ),
  .r_icb_cmd_excl                 (mst_grp_3_ro_icb_cmd_excl                ),
  .r_icb_cmd_xlen                 (mst_grp_3_ro_icb_cmd_xlen     [   7:   0]),
  .r_icb_cmd_xburst               (mst_grp_3_ro_icb_cmd_xburst   [   1:   0]),
  .r_icb_cmd_modes                (mst_grp_3_ro_icb_cmd_modes    [   1:   0]),
  .r_icb_cmd_dmode                (mst_grp_3_ro_icb_cmd_dmode               ),
  .r_icb_cmd_attri                (mst_grp_3_ro_icb_cmd_attri    [   2:   0]),
  .r_icb_cmd_beat                 (mst_grp_3_ro_icb_cmd_beat     [   1:   0]),
  .r_icb_cmd_usr                  (mst_grp_3_ro_icb_cmd_usr      [   2:   0]),
  .r_icb_rsp_ready                (mst_grp_3_ro_icb_rsp_ready               ),
  .r_icb_rsp_valid                (mst_grp_3_ro_icb_rsp_valid               ),
  .r_icb_rsp_err                  (mst_grp_3_ro_icb_rsp_err                 ),
  .r_icb_rsp_excl_ok              (mst_grp_3_ro_icb_rsp_excl_ok             ),
  .r_icb_rsp_rdata                (mst_grp_3_ro_icb_rsp_rdata    [  63:   0]),
  .r_icb_rsp_usr                  (mst_grp_3_ro_icb_rsp_usr      [   2:   0]),
      .w_icb_cmd_valid                (mst_grp_3_wo_icb_cmd_valid               ),
  .w_icb_cmd_ready                (mst_grp_3_wo_icb_cmd_ready               ),
  .w_icb_cmd_sel                  (mst_grp_3_wo_icb_cmd_sel                 ),
  .w_icb_cmd_read                 (mst_grp_3_wo_icb_cmd_read                ),
  .w_icb_cmd_addr                 (mst_grp_3_wo_icb_cmd_addr     [  31:   0]),
  .w_icb_cmd_wdata                (mst_grp_3_wo_icb_cmd_wdata    [  63:   0]),
  .w_icb_cmd_wmask                (mst_grp_3_wo_icb_cmd_wmask    [   7:   0]),
  .w_icb_cmd_size                 (mst_grp_3_wo_icb_cmd_size     [   2:   0]),
  .w_icb_cmd_lock                 (mst_grp_3_wo_icb_cmd_lock                ),
  .w_icb_cmd_excl                 (mst_grp_3_wo_icb_cmd_excl                ),
  .w_icb_cmd_xlen                 (mst_grp_3_wo_icb_cmd_xlen     [   7:   0]),
  .w_icb_cmd_xburst               (mst_grp_3_wo_icb_cmd_xburst   [   1:   0]),
  .w_icb_cmd_modes                (mst_grp_3_wo_icb_cmd_modes    [   1:   0]),
  .w_icb_cmd_dmode                (mst_grp_3_wo_icb_cmd_dmode               ),
  .w_icb_cmd_attri                (mst_grp_3_wo_icb_cmd_attri    [   2:   0]),
  .w_icb_cmd_beat                 (mst_grp_3_wo_icb_cmd_beat     [   1:   0]),
  .w_icb_cmd_usr                  (mst_grp_3_wo_icb_cmd_usr      [   2:   0]),
  .w_icb_rsp_ready                (mst_grp_3_wo_icb_rsp_ready               ),
  .w_icb_rsp_valid                (mst_grp_3_wo_icb_rsp_valid               ),
  .w_icb_rsp_err                  (mst_grp_3_wo_icb_rsp_err                 ),
  .w_icb_rsp_excl_ok              (mst_grp_3_wo_icb_rsp_excl_ok             ),
  .w_icb_rsp_rdata                (mst_grp_3_wo_icb_rsp_rdata    [  63:   0]),
  .w_icb_rsp_usr                  (mst_grp_3_wo_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
      wire                mst_grp_5_ro_icb_cmd_valid    ;
  wire                mst_grp_5_ro_icb_cmd_ready    ;
  wire                mst_grp_5_ro_icb_cmd_sel      ;
  wire                mst_grp_5_ro_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_5_ro_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_5_ro_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_5_ro_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_5_ro_icb_cmd_size     ;
  wire                mst_grp_5_ro_icb_cmd_lock     ;
  wire                mst_grp_5_ro_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_5_ro_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_5_ro_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_5_ro_icb_cmd_modes    ;
  wire                mst_grp_5_ro_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_5_ro_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_5_ro_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_5_ro_icb_cmd_usr      ;
  wire                mst_grp_5_ro_icb_rsp_ready    ;
  wire                mst_grp_5_ro_icb_rsp_valid    ;
  wire                mst_grp_5_ro_icb_rsp_err      ;
  wire                mst_grp_5_ro_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_5_ro_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_5_ro_icb_rsp_usr      ;
      wire                mst_grp_5_wo_icb_cmd_valid    ;
  wire                mst_grp_5_wo_icb_cmd_ready    ;
  wire                mst_grp_5_wo_icb_cmd_sel      ;
  wire                mst_grp_5_wo_icb_cmd_read     ;
  wire    [  31:   0] mst_grp_5_wo_icb_cmd_addr     ;
  wire    [  63:   0] mst_grp_5_wo_icb_cmd_wdata    ;
  wire    [   7:   0] mst_grp_5_wo_icb_cmd_wmask    ;
  wire    [   2:   0] mst_grp_5_wo_icb_cmd_size     ;
  wire                mst_grp_5_wo_icb_cmd_lock     ;
  wire                mst_grp_5_wo_icb_cmd_excl     ;
  wire    [   7:   0] mst_grp_5_wo_icb_cmd_xlen     ;
  wire    [   1:   0] mst_grp_5_wo_icb_cmd_xburst   ;
  wire    [   1:   0] mst_grp_5_wo_icb_cmd_modes    ;
  wire                mst_grp_5_wo_icb_cmd_dmode    ;
  wire    [   2:   0] mst_grp_5_wo_icb_cmd_attri    ;
  wire    [   1:   0] mst_grp_5_wo_icb_cmd_beat     ;
  wire    [   2:   0] mst_grp_5_wo_icb_cmd_usr      ;
  wire                mst_grp_5_wo_icb_rsp_ready    ;
  wire                mst_grp_5_wo_icb_rsp_valid    ;
  wire                mst_grp_5_wo_icb_rsp_err      ;
  wire                mst_grp_5_wo_icb_rsp_excl_ok  ;
  wire    [  63:   0] mst_grp_5_wo_icb_rsp_rdata    ;
  wire    [   2:   0] mst_grp_5_wo_icb_rsp_usr      ;
  e603_subsys_gnrl_ficb_rw_splt # (
      .ALLOW_DIFF   (0),
      .AW           (32),
      .DW           (64),
      .OUTS_FIFO_DP (64),
      .CMD_UW       (3),
      .RSP_UW       (3) 
   ) u_xbar_mg5_rw_splt(
      .icb_cmd_valid                  (mst_grp_5_icb_cmd_valid                  ),
  .icb_cmd_ready                  (mst_grp_5_icb_cmd_ready                  ),
  .icb_cmd_sel                    (mst_grp_5_icb_cmd_sel                    ),
  .icb_cmd_read                   (mst_grp_5_icb_cmd_read                   ),
  .icb_cmd_addr                   (mst_grp_5_icb_cmd_addr        [  31:   0]),
  .icb_cmd_wdata                  (mst_grp_5_icb_cmd_wdata       [  63:   0]),
  .icb_cmd_wmask                  (mst_grp_5_icb_cmd_wmask       [   7:   0]),
  .icb_cmd_size                   (mst_grp_5_icb_cmd_size        [   2:   0]),
  .icb_cmd_lock                   (mst_grp_5_icb_cmd_lock                   ),
  .icb_cmd_excl                   (mst_grp_5_icb_cmd_excl                   ),
  .icb_cmd_xlen                   (mst_grp_5_icb_cmd_xlen        [   7:   0]),
  .icb_cmd_xburst                 (mst_grp_5_icb_cmd_xburst      [   1:   0]),
  .icb_cmd_modes                  (mst_grp_5_icb_cmd_modes       [   1:   0]),
  .icb_cmd_dmode                  (mst_grp_5_icb_cmd_dmode                  ),
  .icb_cmd_attri                  (mst_grp_5_icb_cmd_attri       [   2:   0]),
  .icb_cmd_beat                   (mst_grp_5_icb_cmd_beat        [   1:   0]),
  .icb_cmd_usr                    (mst_grp_5_icb_cmd_usr         [   2:   0]),
  .icb_rsp_ready                  (mst_grp_5_icb_rsp_ready                  ),
  .icb_rsp_valid                  (mst_grp_5_icb_rsp_valid                  ),
  .icb_rsp_err                    (mst_grp_5_icb_rsp_err                    ),
  .icb_rsp_excl_ok                (mst_grp_5_icb_rsp_excl_ok                ),
  .icb_rsp_rdata                  (mst_grp_5_icb_rsp_rdata       [  63:   0]),
  .icb_rsp_usr                    (mst_grp_5_icb_rsp_usr         [   2:   0]),
      .r_icb_cmd_valid                (mst_grp_5_ro_icb_cmd_valid               ),
  .r_icb_cmd_ready                (mst_grp_5_ro_icb_cmd_ready               ),
  .r_icb_cmd_sel                  (mst_grp_5_ro_icb_cmd_sel                 ),
  .r_icb_cmd_read                 (mst_grp_5_ro_icb_cmd_read                ),
  .r_icb_cmd_addr                 (mst_grp_5_ro_icb_cmd_addr     [  31:   0]),
  .r_icb_cmd_wdata                (mst_grp_5_ro_icb_cmd_wdata    [  63:   0]),
  .r_icb_cmd_wmask                (mst_grp_5_ro_icb_cmd_wmask    [   7:   0]),
  .r_icb_cmd_size                 (mst_grp_5_ro_icb_cmd_size     [   2:   0]),
  .r_icb_cmd_lock                 (mst_grp_5_ro_icb_cmd_lock                ),
  .r_icb_cmd_excl                 (mst_grp_5_ro_icb_cmd_excl                ),
  .r_icb_cmd_xlen                 (mst_grp_5_ro_icb_cmd_xlen     [   7:   0]),
  .r_icb_cmd_xburst               (mst_grp_5_ro_icb_cmd_xburst   [   1:   0]),
  .r_icb_cmd_modes                (mst_grp_5_ro_icb_cmd_modes    [   1:   0]),
  .r_icb_cmd_dmode                (mst_grp_5_ro_icb_cmd_dmode               ),
  .r_icb_cmd_attri                (mst_grp_5_ro_icb_cmd_attri    [   2:   0]),
  .r_icb_cmd_beat                 (mst_grp_5_ro_icb_cmd_beat     [   1:   0]),
  .r_icb_cmd_usr                  (mst_grp_5_ro_icb_cmd_usr      [   2:   0]),
  .r_icb_rsp_ready                (mst_grp_5_ro_icb_rsp_ready               ),
  .r_icb_rsp_valid                (mst_grp_5_ro_icb_rsp_valid               ),
  .r_icb_rsp_err                  (mst_grp_5_ro_icb_rsp_err                 ),
  .r_icb_rsp_excl_ok              (mst_grp_5_ro_icb_rsp_excl_ok             ),
  .r_icb_rsp_rdata                (mst_grp_5_ro_icb_rsp_rdata    [  63:   0]),
  .r_icb_rsp_usr                  (mst_grp_5_ro_icb_rsp_usr      [   2:   0]),
      .w_icb_cmd_valid                (mst_grp_5_wo_icb_cmd_valid               ),
  .w_icb_cmd_ready                (mst_grp_5_wo_icb_cmd_ready               ),
  .w_icb_cmd_sel                  (mst_grp_5_wo_icb_cmd_sel                 ),
  .w_icb_cmd_read                 (mst_grp_5_wo_icb_cmd_read                ),
  .w_icb_cmd_addr                 (mst_grp_5_wo_icb_cmd_addr     [  31:   0]),
  .w_icb_cmd_wdata                (mst_grp_5_wo_icb_cmd_wdata    [  63:   0]),
  .w_icb_cmd_wmask                (mst_grp_5_wo_icb_cmd_wmask    [   7:   0]),
  .w_icb_cmd_size                 (mst_grp_5_wo_icb_cmd_size     [   2:   0]),
  .w_icb_cmd_lock                 (mst_grp_5_wo_icb_cmd_lock                ),
  .w_icb_cmd_excl                 (mst_grp_5_wo_icb_cmd_excl                ),
  .w_icb_cmd_xlen                 (mst_grp_5_wo_icb_cmd_xlen     [   7:   0]),
  .w_icb_cmd_xburst               (mst_grp_5_wo_icb_cmd_xburst   [   1:   0]),
  .w_icb_cmd_modes                (mst_grp_5_wo_icb_cmd_modes    [   1:   0]),
  .w_icb_cmd_dmode                (mst_grp_5_wo_icb_cmd_dmode               ),
  .w_icb_cmd_attri                (mst_grp_5_wo_icb_cmd_attri    [   2:   0]),
  .w_icb_cmd_beat                 (mst_grp_5_wo_icb_cmd_beat     [   1:   0]),
  .w_icb_cmd_usr                  (mst_grp_5_wo_icb_cmd_usr      [   2:   0]),
  .w_icb_rsp_ready                (mst_grp_5_wo_icb_rsp_ready               ),
  .w_icb_rsp_valid                (mst_grp_5_wo_icb_rsp_valid               ),
  .w_icb_rsp_err                  (mst_grp_5_wo_icb_rsp_err                 ),
  .w_icb_rsp_excl_ok              (mst_grp_5_wo_icb_rsp_excl_ok             ),
  .w_icb_rsp_rdata                (mst_grp_5_wo_icb_rsp_rdata    [  63:   0]),
  .w_icb_rsp_usr                  (mst_grp_5_wo_icb_rsp_usr      [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst0_ro_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (128  ),
      .SPLT_FIFO_OUTS_CNT_W(8),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg0_ro_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_0_ro_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_0_ro_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_0_ro_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_0_ro_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_0_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_0_ro_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_0_ro_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_0_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_0_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_0_ro_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_0_ro_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_0_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_0_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_0_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_0_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_0_ro_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_0_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_0_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_0_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_0_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_0_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_0_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_0_ro_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg0_ro_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg0_ro_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg0_ro_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg0_ro_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg0_ro_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg0_ro_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg0_ro_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg0_ro_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg0_ro_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg0_ro_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg0_ro_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg0_ro_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg0_ro_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg0_ro_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg0_ro_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg0_ro_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg0_ro_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg0_ro_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg0_ro_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg0_ro_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg0_ro_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg0_ro_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg0_ro_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg0_ro_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg0_ro_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg0_ro_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg0_ro_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg0_ro_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg0_ro_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg0_ro_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg0_ro_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg0_ro_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg0_ro_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg0_ro_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg0_ro_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg0_ro_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg0_ro_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg0_ro_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg0_ro_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg0_ro_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg0_ro_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg0_ro_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg0_ro_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg0_ro_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg0_ro_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg0_ro_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg0_ro_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg0_ro_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg0_ro_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg0_ro_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg0_ro_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg0_ro_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg0_ro_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg0_ro_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg0_ro_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg0_ro_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg0_ro_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg0_ro_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg0_ro_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg0_ro_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg0_ro_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg0_ro_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg0_ro_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg0_ro_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg0_ro_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg0_ro_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg0_ro_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg0_ro_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg0_ro_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg0_ro_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg0_ro_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg0_ro_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg0_ro_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg0_ro_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg0_ro_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg0_ro_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg0_ro_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg0_ro_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg0_ro_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg0_ro_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg0_ro_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg0_ro_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg0_ro_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg0_ro_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg0_ro_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg0_ro_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg0_ro_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg0_ro_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg0_ro_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg0_ro_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg0_ro_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg0_ro_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg0_ro_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg0_ro_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg0_ro_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg0_ro_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg0_ro_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg0_ro_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg0_ro_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg0_ro_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg0_ro_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg0_ro_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg0_ro_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg0_ro_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg0_ro_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg0_ro_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg0_ro_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg0_ro_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg0_ro_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg0_ro_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg0_ro_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg0_ro_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg0_ro_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg0_ro_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg0_ro_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg0_ro_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg0_ro_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg0_ro_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg0_ro_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg0_ro_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg0_ro_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg0_ro_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg0_ro_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg0_ro_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg0_ro_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg0_ro_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg0_ro_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg0_ro_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg0_ro_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg0_ro_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg0_ro_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg0_ro_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg0_ro_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg0_ro_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg0_ro_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg0_ro_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg0_ro_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg0_ro_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg0_ro_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg0_ro_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg0_ro_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg0_ro_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg0_ro_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg0_ro_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg0_ro_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg0_ro_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg0_ro_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg0_ro_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg0_ro_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg0_ro_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg0_ro_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg0_ro_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg0_ro_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg0_ro_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst1_ro_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg1_ro_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_1_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (mst_grp_1_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (mst_grp_1_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (mst_grp_1_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (mst_grp_1_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_1_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_1_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_1_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_1_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (mst_grp_1_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (mst_grp_1_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_1_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_1_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_1_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (mst_grp_1_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_1_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_1_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_1_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (mst_grp_1_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (mst_grp_1_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (mst_grp_1_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (mst_grp_1_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_1_icb_rsp_usr         [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg1_ro_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg1_ro_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg1_ro_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg1_ro_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg1_ro_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg1_ro_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg1_ro_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg1_ro_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg1_ro_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg1_ro_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg1_ro_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg1_ro_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg1_ro_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg1_ro_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg1_ro_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg1_ro_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg1_ro_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg1_ro_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg1_ro_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg1_ro_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg1_ro_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg1_ro_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg1_ro_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg1_ro_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg1_ro_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg1_ro_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg1_ro_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg1_ro_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg1_ro_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg1_ro_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg1_ro_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg1_ro_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg1_ro_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg1_ro_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg1_ro_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg1_ro_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg1_ro_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg1_ro_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg1_ro_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg1_ro_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg1_ro_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg1_ro_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg1_ro_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg1_ro_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg1_ro_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg1_ro_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg1_ro_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg1_ro_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg1_ro_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg1_ro_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg1_ro_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg1_ro_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg1_ro_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg1_ro_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg1_ro_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg1_ro_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg1_ro_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg1_ro_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg1_ro_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg1_ro_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg1_ro_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg1_ro_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg1_ro_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg1_ro_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg1_ro_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg1_ro_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg1_ro_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg1_ro_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg1_ro_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg1_ro_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg1_ro_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg1_ro_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg1_ro_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg1_ro_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg1_ro_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg1_ro_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg1_ro_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg1_ro_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg1_ro_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg1_ro_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg1_ro_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg1_ro_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg1_ro_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg1_ro_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg1_ro_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg1_ro_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg1_ro_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg1_ro_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg1_ro_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg1_ro_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg1_ro_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg1_ro_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg1_ro_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg1_ro_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg1_ro_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg1_ro_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg1_ro_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg1_ro_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg1_ro_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg1_ro_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg1_ro_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg1_ro_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg1_ro_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg1_ro_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg1_ro_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg1_ro_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg1_ro_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg1_ro_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg1_ro_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg1_ro_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg1_ro_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg1_ro_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg1_ro_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg1_ro_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg1_ro_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg1_ro_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg1_ro_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg1_ro_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg1_ro_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg1_ro_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg1_ro_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg1_ro_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg1_ro_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg1_ro_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg1_ro_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg1_ro_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg1_ro_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg1_ro_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg1_ro_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg1_ro_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg1_ro_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg1_ro_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg1_ro_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg1_ro_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg1_ro_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg1_ro_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg1_ro_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg1_ro_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg1_ro_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg1_ro_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg1_ro_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg1_ro_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg1_ro_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg1_ro_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg1_ro_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg1_ro_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg1_ro_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg1_ro_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg1_ro_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg1_ro_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg1_ro_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg1_ro_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg1_ro_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg1_ro_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst3_ro_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg3_ro_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_3_ro_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_3_ro_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_3_ro_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_3_ro_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_3_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_3_ro_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_3_ro_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_3_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_3_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_3_ro_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_3_ro_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_3_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_3_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_3_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_3_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_3_ro_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_3_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_3_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_3_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_3_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_3_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_3_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_3_ro_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg3_ro_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg3_ro_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg3_ro_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg3_ro_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg3_ro_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg3_ro_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg3_ro_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg3_ro_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg3_ro_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg3_ro_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg3_ro_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg3_ro_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg3_ro_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg3_ro_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg3_ro_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg3_ro_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg3_ro_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg3_ro_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg3_ro_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg3_ro_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg3_ro_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg3_ro_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg3_ro_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg3_ro_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg3_ro_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg3_ro_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg3_ro_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg3_ro_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg3_ro_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg3_ro_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg3_ro_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg3_ro_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg3_ro_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg3_ro_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg3_ro_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg3_ro_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg3_ro_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg3_ro_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg3_ro_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg3_ro_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg3_ro_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg3_ro_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg3_ro_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg3_ro_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg3_ro_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg3_ro_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg3_ro_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg3_ro_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg3_ro_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg3_ro_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg3_ro_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg3_ro_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg3_ro_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg3_ro_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg3_ro_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg3_ro_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg3_ro_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg3_ro_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg3_ro_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg3_ro_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg3_ro_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg3_ro_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg3_ro_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg3_ro_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg3_ro_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg3_ro_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg3_ro_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg3_ro_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg3_ro_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg3_ro_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg3_ro_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg3_ro_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg3_ro_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg3_ro_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg3_ro_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg3_ro_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg3_ro_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg3_ro_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg3_ro_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg3_ro_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg3_ro_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg3_ro_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg3_ro_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg3_ro_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg3_ro_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg3_ro_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg3_ro_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg3_ro_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg3_ro_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg3_ro_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg3_ro_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg3_ro_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg3_ro_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg3_ro_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg3_ro_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg3_ro_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg3_ro_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg3_ro_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg3_ro_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg3_ro_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg3_ro_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg3_ro_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg3_ro_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg3_ro_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg3_ro_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg3_ro_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg3_ro_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg3_ro_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg3_ro_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg3_ro_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg3_ro_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg3_ro_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg3_ro_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg3_ro_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg3_ro_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg3_ro_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg3_ro_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg3_ro_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg3_ro_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg3_ro_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg3_ro_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg3_ro_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg3_ro_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg3_ro_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg3_ro_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg3_ro_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg3_ro_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg3_ro_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg3_ro_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg3_ro_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg3_ro_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg3_ro_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg3_ro_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg3_ro_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg3_ro_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg3_ro_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg3_ro_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg3_ro_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg3_ro_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg3_ro_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg3_ro_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg3_ro_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg3_ro_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg3_ro_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg3_ro_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg3_ro_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg3_ro_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg3_ro_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg3_ro_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg3_ro_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg3_ro_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg3_ro_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg3_ro_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg3_ro_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst4_ro_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg4_ro_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_4_ro_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_4_ro_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_4_ro_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_4_ro_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_4_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_4_ro_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_4_ro_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_4_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_4_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_4_ro_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_4_ro_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_4_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_4_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_4_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_4_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_4_ro_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_4_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_4_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_4_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_4_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_4_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_4_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_4_ro_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg4_ro_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg4_ro_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg4_ro_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg4_ro_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg4_ro_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg4_ro_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg4_ro_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg4_ro_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg4_ro_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg4_ro_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg4_ro_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg4_ro_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg4_ro_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg4_ro_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg4_ro_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg4_ro_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg4_ro_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg4_ro_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg4_ro_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg4_ro_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg4_ro_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg4_ro_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg4_ro_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg4_ro_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg4_ro_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg4_ro_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg4_ro_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg4_ro_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg4_ro_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg4_ro_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg4_ro_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg4_ro_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg4_ro_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg4_ro_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg4_ro_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg4_ro_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg4_ro_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg4_ro_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg4_ro_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg4_ro_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg4_ro_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg4_ro_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg4_ro_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg4_ro_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg4_ro_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg4_ro_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg4_ro_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg4_ro_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg4_ro_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg4_ro_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg4_ro_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg4_ro_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg4_ro_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg4_ro_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg4_ro_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg4_ro_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg4_ro_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg4_ro_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg4_ro_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg4_ro_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg4_ro_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg4_ro_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg4_ro_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg4_ro_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg4_ro_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg4_ro_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg4_ro_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg4_ro_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg4_ro_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg4_ro_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg4_ro_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg4_ro_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg4_ro_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg4_ro_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg4_ro_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg4_ro_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg4_ro_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg4_ro_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg4_ro_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg4_ro_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg4_ro_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg4_ro_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg4_ro_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg4_ro_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg4_ro_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg4_ro_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg4_ro_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg4_ro_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg4_ro_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg4_ro_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg4_ro_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg4_ro_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg4_ro_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg4_ro_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg4_ro_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg4_ro_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg4_ro_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg4_ro_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg4_ro_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg4_ro_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg4_ro_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg4_ro_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg4_ro_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg4_ro_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg4_ro_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg4_ro_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg4_ro_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg4_ro_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg4_ro_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg4_ro_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg4_ro_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg4_ro_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg4_ro_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg4_ro_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg4_ro_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg4_ro_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg4_ro_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg4_ro_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg4_ro_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg4_ro_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg4_ro_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg4_ro_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg4_ro_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg4_ro_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg4_ro_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg4_ro_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg4_ro_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg4_ro_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg4_ro_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg4_ro_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg4_ro_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg4_ro_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg4_ro_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg4_ro_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg4_ro_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg4_ro_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg4_ro_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg4_ro_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg4_ro_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg4_ro_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg4_ro_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg4_ro_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg4_ro_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg4_ro_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg4_ro_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg4_ro_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg4_ro_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg4_ro_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg4_ro_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg4_ro_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg4_ro_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg4_ro_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg4_ro_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg4_ro_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst5_ro_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg5_ro_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_5_ro_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_5_ro_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_5_ro_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_5_ro_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_5_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_5_ro_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_5_ro_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_5_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_5_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_5_ro_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_5_ro_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_5_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_5_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_5_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_5_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_5_ro_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_5_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_5_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_5_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_5_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_5_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_5_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_5_ro_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg5_ro_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg5_ro_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg5_ro_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg5_ro_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg5_ro_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg5_ro_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg5_ro_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg5_ro_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg5_ro_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg5_ro_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg5_ro_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg5_ro_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg5_ro_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg5_ro_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg5_ro_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg5_ro_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg5_ro_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg5_ro_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg5_ro_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg5_ro_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg5_ro_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg5_ro_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg5_ro_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg5_ro_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg5_ro_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg5_ro_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg5_ro_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg5_ro_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg5_ro_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg5_ro_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg5_ro_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg5_ro_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg5_ro_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg5_ro_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg5_ro_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg5_ro_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg5_ro_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg5_ro_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg5_ro_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg5_ro_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg5_ro_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg5_ro_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg5_ro_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg5_ro_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg5_ro_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg5_ro_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg5_ro_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg5_ro_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg5_ro_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg5_ro_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg5_ro_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg5_ro_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg5_ro_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg5_ro_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg5_ro_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg5_ro_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg5_ro_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg5_ro_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg5_ro_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg5_ro_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg5_ro_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg5_ro_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg5_ro_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg5_ro_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg5_ro_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg5_ro_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg5_ro_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg5_ro_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg5_ro_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg5_ro_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg5_ro_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg5_ro_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg5_ro_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg5_ro_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg5_ro_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg5_ro_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg5_ro_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg5_ro_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg5_ro_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg5_ro_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg5_ro_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg5_ro_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg5_ro_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg5_ro_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg5_ro_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg5_ro_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg5_ro_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg5_ro_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg5_ro_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg5_ro_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg5_ro_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg5_ro_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg5_ro_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg5_ro_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg5_ro_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg5_ro_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg5_ro_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg5_ro_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg5_ro_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg5_ro_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg5_ro_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg5_ro_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg5_ro_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg5_ro_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg5_ro_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg5_ro_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg5_ro_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg5_ro_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg5_ro_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg5_ro_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg5_ro_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg5_ro_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg5_ro_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg5_ro_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg5_ro_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg5_ro_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg5_ro_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg5_ro_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg5_ro_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg5_ro_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg5_ro_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg5_ro_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg5_ro_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg5_ro_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg5_ro_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg5_ro_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg5_ro_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg5_ro_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg5_ro_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg5_ro_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg5_ro_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg5_ro_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg5_ro_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg5_ro_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg5_ro_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg5_ro_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg5_ro_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg5_ro_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg5_ro_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg5_ro_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg5_ro_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg5_ro_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg5_ro_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg5_ro_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg5_ro_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg5_ro_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg5_ro_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg5_ro_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg5_ro_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg5_ro_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg5_ro_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg5_ro_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg5_ro_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg5_ro_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst6_ro_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg6_ro_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_6_ro_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_6_ro_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_6_ro_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_6_ro_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_6_ro_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_6_ro_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_6_ro_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_6_ro_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_6_ro_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_6_ro_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_6_ro_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_6_ro_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_6_ro_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_6_ro_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_6_ro_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_6_ro_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_6_ro_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_6_ro_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_6_ro_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_6_ro_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_6_ro_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_6_ro_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_6_ro_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg6_ro_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg6_ro_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg6_ro_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg6_ro_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg6_ro_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg6_ro_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg6_ro_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg6_ro_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg6_ro_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg6_ro_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg6_ro_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg6_ro_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg6_ro_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg6_ro_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg6_ro_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg6_ro_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg6_ro_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg6_ro_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg6_ro_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg6_ro_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg6_ro_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg6_ro_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg6_ro_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg6_ro_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg6_ro_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg6_ro_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg6_ro_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg6_ro_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg6_ro_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg6_ro_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg6_ro_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg6_ro_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg6_ro_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg6_ro_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg6_ro_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg6_ro_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg6_ro_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg6_ro_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg6_ro_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg6_ro_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg6_ro_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg6_ro_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg6_ro_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg6_ro_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg6_ro_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg6_ro_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg6_ro_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg6_ro_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg6_ro_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg6_ro_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg6_ro_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg6_ro_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg6_ro_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg6_ro_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg6_ro_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg6_ro_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg6_ro_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg6_ro_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg6_ro_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg6_ro_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg6_ro_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg6_ro_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg6_ro_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg6_ro_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg6_ro_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg6_ro_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg6_ro_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg6_ro_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg6_ro_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg6_ro_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg6_ro_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg6_ro_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg6_ro_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg6_ro_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg6_ro_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg6_ro_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg6_ro_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg6_ro_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg6_ro_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg6_ro_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg6_ro_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg6_ro_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg6_ro_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg6_ro_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg6_ro_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg6_ro_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg6_ro_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg6_ro_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg6_ro_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg6_ro_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg6_ro_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg6_ro_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg6_ro_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg6_ro_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg6_ro_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg6_ro_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg6_ro_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg6_ro_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg6_ro_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg6_ro_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg6_ro_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg6_ro_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg6_ro_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg6_ro_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg6_ro_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg6_ro_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg6_ro_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg6_ro_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg6_ro_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg6_ro_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg6_ro_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg6_ro_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg6_ro_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg6_ro_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg6_ro_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg6_ro_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg6_ro_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg6_ro_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg6_ro_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg6_ro_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg6_ro_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg6_ro_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg6_ro_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg6_ro_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg6_ro_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg6_ro_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg6_ro_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg6_ro_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg6_ro_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg6_ro_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg6_ro_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg6_ro_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg6_ro_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg6_ro_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg6_ro_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg6_ro_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg6_ro_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg6_ro_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg6_ro_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg6_ro_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg6_ro_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg6_ro_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg6_ro_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg6_ro_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg6_ro_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg6_ro_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg6_ro_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg6_ro_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg6_ro_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg6_ro_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg6_ro_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg6_ro_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg6_ro_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg6_ro_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst0_wo_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (128  ),
      .SPLT_FIFO_OUTS_CNT_W(8),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg0_wo_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_0_wo_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_0_wo_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_0_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_0_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_0_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_0_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_0_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_0_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_0_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_0_wo_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_0_wo_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_0_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_0_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_0_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_0_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_0_wo_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_0_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_0_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_0_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_0_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_0_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_0_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_0_wo_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg0_wo_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg0_wo_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg0_wo_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg0_wo_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg0_wo_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg0_wo_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg0_wo_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg0_wo_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg0_wo_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg0_wo_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg0_wo_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg0_wo_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg0_wo_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg0_wo_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg0_wo_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg0_wo_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg0_wo_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg0_wo_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg0_wo_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg0_wo_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg0_wo_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg0_wo_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg0_wo_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg0_wo_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg0_wo_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg0_wo_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg0_wo_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg0_wo_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg0_wo_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg0_wo_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg0_wo_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg0_wo_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg0_wo_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg0_wo_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg0_wo_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg0_wo_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg0_wo_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg0_wo_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg0_wo_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg0_wo_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg0_wo_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg0_wo_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg0_wo_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg0_wo_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg0_wo_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg0_wo_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg0_wo_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg0_wo_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg0_wo_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg0_wo_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg0_wo_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg0_wo_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg0_wo_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg0_wo_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg0_wo_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg0_wo_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg0_wo_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg0_wo_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg0_wo_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg0_wo_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg0_wo_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg0_wo_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg0_wo_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg0_wo_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg0_wo_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg0_wo_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg0_wo_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg0_wo_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg0_wo_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg0_wo_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg0_wo_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg0_wo_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg0_wo_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg0_wo_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg0_wo_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg0_wo_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg0_wo_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg0_wo_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg0_wo_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg0_wo_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg0_wo_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg0_wo_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg0_wo_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg0_wo_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg0_wo_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg0_wo_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg0_wo_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg0_wo_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg0_wo_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg0_wo_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg0_wo_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg0_wo_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg0_wo_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg0_wo_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg0_wo_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg0_wo_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg0_wo_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg0_wo_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg0_wo_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg0_wo_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg0_wo_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg0_wo_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg0_wo_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg0_wo_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg0_wo_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg0_wo_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg0_wo_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg0_wo_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg0_wo_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg0_wo_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg0_wo_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg0_wo_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg0_wo_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg0_wo_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg0_wo_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg0_wo_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg0_wo_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg0_wo_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg0_wo_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg0_wo_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg0_wo_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg0_wo_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg0_wo_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg0_wo_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg0_wo_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg0_wo_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg0_wo_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg0_wo_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg0_wo_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg0_wo_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg0_wo_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg0_wo_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg0_wo_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg0_wo_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg0_wo_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg0_wo_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg0_wo_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg0_wo_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg0_wo_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg0_wo_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg0_wo_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg0_wo_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg0_wo_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg0_wo_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg0_wo_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg0_wo_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg0_wo_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg0_wo_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg0_wo_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg0_wo_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg0_wo_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg0_wo_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg0_wo_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg0_wo_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst2_wo_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg2_wo_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_2_icb_cmd_valid                  ),
  .i_icb_cmd_ready                (mst_grp_2_icb_cmd_ready                  ),
  .i_icb_cmd_sel                  (mst_grp_2_icb_cmd_sel                    ),
  .i_icb_cmd_read                 (mst_grp_2_icb_cmd_read                   ),
  .i_icb_cmd_addr                 (mst_grp_2_icb_cmd_addr        [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_2_icb_cmd_wdata       [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_2_icb_cmd_wmask       [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_2_icb_cmd_size        [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_2_icb_cmd_lock                   ),
  .i_icb_cmd_excl                 (mst_grp_2_icb_cmd_excl                   ),
  .i_icb_cmd_xlen                 (mst_grp_2_icb_cmd_xlen        [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_2_icb_cmd_xburst      [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_2_icb_cmd_modes       [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_2_icb_cmd_dmode                  ),
  .i_icb_cmd_attri                (mst_grp_2_icb_cmd_attri       [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_2_icb_cmd_beat        [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_2_icb_cmd_usr         [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_2_icb_rsp_ready                  ),
  .i_icb_rsp_valid                (mst_grp_2_icb_rsp_valid                  ),
  .i_icb_rsp_err                  (mst_grp_2_icb_rsp_err                    ),
  .i_icb_rsp_excl_ok              (mst_grp_2_icb_rsp_excl_ok                ),
  .i_icb_rsp_rdata                (mst_grp_2_icb_rsp_rdata       [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_2_icb_rsp_usr         [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg2_wo_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg2_wo_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg2_wo_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg2_wo_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg2_wo_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg2_wo_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg2_wo_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg2_wo_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg2_wo_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg2_wo_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg2_wo_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg2_wo_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg2_wo_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg2_wo_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg2_wo_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg2_wo_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg2_wo_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg2_wo_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg2_wo_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg2_wo_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg2_wo_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg2_wo_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg2_wo_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg2_wo_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg2_wo_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg2_wo_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg2_wo_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg2_wo_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg2_wo_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg2_wo_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg2_wo_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg2_wo_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg2_wo_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg2_wo_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg2_wo_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg2_wo_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg2_wo_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg2_wo_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg2_wo_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg2_wo_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg2_wo_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg2_wo_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg2_wo_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg2_wo_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg2_wo_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg2_wo_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg2_wo_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg2_wo_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg2_wo_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg2_wo_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg2_wo_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg2_wo_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg2_wo_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg2_wo_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg2_wo_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg2_wo_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg2_wo_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg2_wo_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg2_wo_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg2_wo_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg2_wo_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg2_wo_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg2_wo_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg2_wo_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg2_wo_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg2_wo_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg2_wo_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg2_wo_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg2_wo_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg2_wo_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg2_wo_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg2_wo_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg2_wo_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg2_wo_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg2_wo_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg2_wo_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg2_wo_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg2_wo_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg2_wo_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg2_wo_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg2_wo_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg2_wo_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg2_wo_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg2_wo_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg2_wo_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg2_wo_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg2_wo_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg2_wo_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg2_wo_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg2_wo_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg2_wo_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg2_wo_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg2_wo_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg2_wo_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg2_wo_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg2_wo_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg2_wo_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg2_wo_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg2_wo_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg2_wo_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg2_wo_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg2_wo_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg2_wo_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg2_wo_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg2_wo_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg2_wo_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg2_wo_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg2_wo_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg2_wo_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg2_wo_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg2_wo_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg2_wo_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg2_wo_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg2_wo_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg2_wo_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg2_wo_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg2_wo_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg2_wo_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg2_wo_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg2_wo_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg2_wo_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg2_wo_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg2_wo_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg2_wo_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg2_wo_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg2_wo_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg2_wo_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg2_wo_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg2_wo_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg2_wo_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg2_wo_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg2_wo_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg2_wo_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg2_wo_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg2_wo_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg2_wo_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg2_wo_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg2_wo_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg2_wo_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg2_wo_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg2_wo_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg2_wo_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg2_wo_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg2_wo_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg2_wo_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg2_wo_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg2_wo_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg2_wo_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg2_wo_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg2_wo_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg2_wo_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg2_wo_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg2_wo_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg2_wo_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst3_wo_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg3_wo_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_3_wo_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_3_wo_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_3_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_3_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_3_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_3_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_3_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_3_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_3_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_3_wo_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_3_wo_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_3_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_3_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_3_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_3_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_3_wo_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_3_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_3_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_3_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_3_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_3_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_3_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_3_wo_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg3_wo_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg3_wo_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg3_wo_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg3_wo_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg3_wo_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg3_wo_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg3_wo_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg3_wo_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg3_wo_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg3_wo_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg3_wo_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg3_wo_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg3_wo_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg3_wo_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg3_wo_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg3_wo_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg3_wo_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg3_wo_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg3_wo_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg3_wo_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg3_wo_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg3_wo_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg3_wo_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg3_wo_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg3_wo_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg3_wo_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg3_wo_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg3_wo_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg3_wo_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg3_wo_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg3_wo_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg3_wo_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg3_wo_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg3_wo_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg3_wo_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg3_wo_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg3_wo_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg3_wo_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg3_wo_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg3_wo_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg3_wo_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg3_wo_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg3_wo_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg3_wo_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg3_wo_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg3_wo_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg3_wo_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg3_wo_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg3_wo_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg3_wo_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg3_wo_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg3_wo_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg3_wo_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg3_wo_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg3_wo_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg3_wo_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg3_wo_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg3_wo_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg3_wo_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg3_wo_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg3_wo_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg3_wo_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg3_wo_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg3_wo_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg3_wo_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg3_wo_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg3_wo_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg3_wo_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg3_wo_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg3_wo_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg3_wo_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg3_wo_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg3_wo_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg3_wo_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg3_wo_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg3_wo_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg3_wo_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg3_wo_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg3_wo_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg3_wo_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg3_wo_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg3_wo_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg3_wo_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg3_wo_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg3_wo_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg3_wo_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg3_wo_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg3_wo_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg3_wo_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg3_wo_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg3_wo_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg3_wo_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg3_wo_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg3_wo_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg3_wo_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg3_wo_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg3_wo_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg3_wo_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg3_wo_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg3_wo_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg3_wo_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg3_wo_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg3_wo_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg3_wo_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg3_wo_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg3_wo_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg3_wo_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg3_wo_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg3_wo_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg3_wo_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg3_wo_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg3_wo_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg3_wo_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg3_wo_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg3_wo_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg3_wo_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg3_wo_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg3_wo_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg3_wo_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg3_wo_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg3_wo_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg3_wo_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg3_wo_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg3_wo_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg3_wo_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg3_wo_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg3_wo_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg3_wo_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg3_wo_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg3_wo_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg3_wo_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg3_wo_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg3_wo_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg3_wo_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg3_wo_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg3_wo_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg3_wo_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg3_wo_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg3_wo_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg3_wo_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg3_wo_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg3_wo_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg3_wo_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg3_wo_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg3_wo_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg3_wo_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg3_wo_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg3_wo_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg3_wo_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg3_wo_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg3_wo_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg3_wo_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg3_wo_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg3_wo_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst4_wo_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg4_wo_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_4_wo_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_4_wo_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_4_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_4_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_4_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_4_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_4_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_4_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_4_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_4_wo_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_4_wo_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_4_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_4_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_4_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_4_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_4_wo_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_4_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_4_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_4_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_4_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_4_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_4_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_4_wo_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg4_wo_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg4_wo_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg4_wo_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg4_wo_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg4_wo_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg4_wo_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg4_wo_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg4_wo_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg4_wo_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg4_wo_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg4_wo_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg4_wo_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg4_wo_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg4_wo_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg4_wo_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg4_wo_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg4_wo_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg4_wo_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg4_wo_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg4_wo_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg4_wo_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg4_wo_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg4_wo_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg4_wo_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg4_wo_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg4_wo_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg4_wo_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg4_wo_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg4_wo_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg4_wo_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg4_wo_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg4_wo_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg4_wo_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg4_wo_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg4_wo_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg4_wo_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg4_wo_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg4_wo_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg4_wo_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg4_wo_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg4_wo_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg4_wo_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg4_wo_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg4_wo_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg4_wo_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg4_wo_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg4_wo_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg4_wo_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg4_wo_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg4_wo_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg4_wo_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg4_wo_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg4_wo_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg4_wo_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg4_wo_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg4_wo_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg4_wo_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg4_wo_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg4_wo_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg4_wo_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg4_wo_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg4_wo_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg4_wo_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg4_wo_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg4_wo_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg4_wo_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg4_wo_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg4_wo_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg4_wo_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg4_wo_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg4_wo_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg4_wo_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg4_wo_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg4_wo_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg4_wo_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg4_wo_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg4_wo_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg4_wo_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg4_wo_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg4_wo_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg4_wo_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg4_wo_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg4_wo_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg4_wo_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg4_wo_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg4_wo_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg4_wo_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg4_wo_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg4_wo_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg4_wo_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg4_wo_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg4_wo_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg4_wo_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg4_wo_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg4_wo_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg4_wo_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg4_wo_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg4_wo_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg4_wo_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg4_wo_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg4_wo_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg4_wo_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg4_wo_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg4_wo_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg4_wo_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg4_wo_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg4_wo_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg4_wo_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg4_wo_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg4_wo_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg4_wo_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg4_wo_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg4_wo_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg4_wo_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg4_wo_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg4_wo_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg4_wo_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg4_wo_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg4_wo_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg4_wo_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg4_wo_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg4_wo_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg4_wo_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg4_wo_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg4_wo_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg4_wo_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg4_wo_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg4_wo_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg4_wo_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg4_wo_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg4_wo_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg4_wo_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg4_wo_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg4_wo_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg4_wo_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg4_wo_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg4_wo_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg4_wo_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg4_wo_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg4_wo_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg4_wo_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg4_wo_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg4_wo_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg4_wo_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg4_wo_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg4_wo_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg4_wo_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg4_wo_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg4_wo_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg4_wo_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg4_wo_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg4_wo_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg4_wo_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg4_wo_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst5_wo_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg5_wo_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_5_wo_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_5_wo_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_5_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_5_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_5_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_5_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_5_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_5_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_5_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_5_wo_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_5_wo_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_5_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_5_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_5_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_5_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_5_wo_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_5_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_5_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_5_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_5_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_5_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_5_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_5_wo_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg5_wo_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg5_wo_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg5_wo_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg5_wo_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg5_wo_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg5_wo_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg5_wo_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg5_wo_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg5_wo_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg5_wo_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg5_wo_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg5_wo_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg5_wo_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg5_wo_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg5_wo_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg5_wo_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg5_wo_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg5_wo_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg5_wo_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg5_wo_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg5_wo_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg5_wo_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg5_wo_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg5_wo_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg5_wo_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg5_wo_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg5_wo_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg5_wo_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg5_wo_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg5_wo_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg5_wo_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg5_wo_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg5_wo_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg5_wo_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg5_wo_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg5_wo_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg5_wo_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg5_wo_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg5_wo_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg5_wo_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg5_wo_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg5_wo_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg5_wo_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg5_wo_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg5_wo_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg5_wo_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg5_wo_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg5_wo_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg5_wo_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg5_wo_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg5_wo_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg5_wo_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg5_wo_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg5_wo_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg5_wo_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg5_wo_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg5_wo_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg5_wo_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg5_wo_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg5_wo_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg5_wo_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg5_wo_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg5_wo_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg5_wo_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg5_wo_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg5_wo_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg5_wo_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg5_wo_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg5_wo_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg5_wo_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg5_wo_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg5_wo_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg5_wo_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg5_wo_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg5_wo_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg5_wo_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg5_wo_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg5_wo_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg5_wo_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg5_wo_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg5_wo_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg5_wo_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg5_wo_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg5_wo_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg5_wo_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg5_wo_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg5_wo_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg5_wo_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg5_wo_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg5_wo_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg5_wo_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg5_wo_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg5_wo_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg5_wo_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg5_wo_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg5_wo_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg5_wo_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg5_wo_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg5_wo_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg5_wo_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg5_wo_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg5_wo_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg5_wo_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg5_wo_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg5_wo_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg5_wo_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg5_wo_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg5_wo_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg5_wo_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg5_wo_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg5_wo_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg5_wo_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg5_wo_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg5_wo_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg5_wo_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg5_wo_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg5_wo_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg5_wo_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg5_wo_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg5_wo_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg5_wo_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg5_wo_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg5_wo_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg5_wo_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg5_wo_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg5_wo_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg5_wo_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg5_wo_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg5_wo_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg5_wo_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg5_wo_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg5_wo_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg5_wo_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg5_wo_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg5_wo_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg5_wo_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg5_wo_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg5_wo_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg5_wo_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg5_wo_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg5_wo_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg5_wo_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg5_wo_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg5_wo_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg5_wo_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg5_wo_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg5_wo_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg5_wo_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg5_wo_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg5_wo_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg5_wo_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg5_wo_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg5_wo_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg5_wo_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
   e603_subsys_xbar_mst6_wo_ficb1ton_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ALLOW_DIFF             (0),
      .ALLOW_0CYCL_RSP        (0),
      .ICB_FIFO_CMD_BYPBUF    (1), 
      .ICB_FIFO_CMD_DP        (1), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .O0_BASE_ADDR       (32'h60000000),
      .O0_BASE_REGION_LSB (16),
      .O1_BASE_ADDR       (32'h68000000),
      .O1_BASE_REGION_LSB (16),
      .O2_BASE_ADDR       (32'h0),
      .O2_BASE_REGION_LSB (12),
      .O3_BASE_ADDR       (32'h20000000),
      .O3_BASE_REGION_LSB (28),
      .O4_BASE_ADDR       (32'h10000000),
      .O4_BASE_REGION_LSB (20),
      .O5_BASE_ADDR       (32'h80000000),
      .O5_BASE_REGION_LSB (31),
      .O6_BASE_ADDR       (0),
      .O6_BASE_REGION_LSB (0),
      .SPLT_FIFO_OUTS_NUM  (64  ),
      .SPLT_FIFO_OUTS_CNT_W(7),
      .SPLT_FIFO_CUT_READY (1) 
   ) u_xbar_mg6_wo_icb1ton(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icb1ton_active (),
      .i_icb_cmd_valid                (mst_grp_6_wo_icb_cmd_valid               ),
  .i_icb_cmd_ready                (mst_grp_6_wo_icb_cmd_ready               ),
  .i_icb_cmd_sel                  (mst_grp_6_wo_icb_cmd_sel                 ),
  .i_icb_cmd_read                 (mst_grp_6_wo_icb_cmd_read                ),
  .i_icb_cmd_addr                 (mst_grp_6_wo_icb_cmd_addr     [  31:   0]),
  .i_icb_cmd_wdata                (mst_grp_6_wo_icb_cmd_wdata    [  63:   0]),
  .i_icb_cmd_wmask                (mst_grp_6_wo_icb_cmd_wmask    [   7:   0]),
  .i_icb_cmd_size                 (mst_grp_6_wo_icb_cmd_size     [   2:   0]),
  .i_icb_cmd_lock                 (mst_grp_6_wo_icb_cmd_lock                ),
  .i_icb_cmd_excl                 (mst_grp_6_wo_icb_cmd_excl                ),
  .i_icb_cmd_xlen                 (mst_grp_6_wo_icb_cmd_xlen     [   7:   0]),
  .i_icb_cmd_xburst               (mst_grp_6_wo_icb_cmd_xburst   [   1:   0]),
  .i_icb_cmd_modes                (mst_grp_6_wo_icb_cmd_modes    [   1:   0]),
  .i_icb_cmd_dmode                (mst_grp_6_wo_icb_cmd_dmode               ),
  .i_icb_cmd_attri                (mst_grp_6_wo_icb_cmd_attri    [   2:   0]),
  .i_icb_cmd_beat                 (mst_grp_6_wo_icb_cmd_beat     [   1:   0]),
  .i_icb_cmd_usr                  (mst_grp_6_wo_icb_cmd_usr      [   2:   0]),
  .i_icb_rsp_ready                (mst_grp_6_wo_icb_rsp_ready               ),
  .i_icb_rsp_valid                (mst_grp_6_wo_icb_rsp_valid               ),
  .i_icb_rsp_err                  (mst_grp_6_wo_icb_rsp_err                 ),
  .i_icb_rsp_excl_ok              (mst_grp_6_wo_icb_rsp_excl_ok             ),
  .i_icb_rsp_rdata                (mst_grp_6_wo_icb_rsp_rdata    [  63:   0]),
  .i_icb_rsp_usr                  (mst_grp_6_wo_icb_rsp_usr      [   2:   0]),
      .o0_icb_enable(1'b1),
      .o0_icb_cmd_valid               (xbar_mg6_wo_to_sg0_cmd_valid             ),
  .o0_icb_cmd_ready               (xbar_mg6_wo_to_sg0_cmd_ready             ),
  .o0_icb_cmd_sel                 (xbar_mg6_wo_to_sg0_cmd_sel               ),
  .o0_icb_cmd_read                (xbar_mg6_wo_to_sg0_cmd_read              ),
  .o0_icb_cmd_addr                (xbar_mg6_wo_to_sg0_cmd_addr   [  31:   0]),
  .o0_icb_cmd_wdata               (xbar_mg6_wo_to_sg0_cmd_wdata  [  63:   0]),
  .o0_icb_cmd_wmask               (xbar_mg6_wo_to_sg0_cmd_wmask  [   7:   0]),
  .o0_icb_cmd_size                (xbar_mg6_wo_to_sg0_cmd_size   [   2:   0]),
  .o0_icb_cmd_lock                (xbar_mg6_wo_to_sg0_cmd_lock              ),
  .o0_icb_cmd_excl                (xbar_mg6_wo_to_sg0_cmd_excl              ),
  .o0_icb_cmd_xlen                (xbar_mg6_wo_to_sg0_cmd_xlen   [   7:   0]),
  .o0_icb_cmd_xburst              (xbar_mg6_wo_to_sg0_cmd_xburst [   1:   0]),
  .o0_icb_cmd_modes               (xbar_mg6_wo_to_sg0_cmd_modes  [   1:   0]),
  .o0_icb_cmd_dmode               (xbar_mg6_wo_to_sg0_cmd_dmode             ),
  .o0_icb_cmd_attri               (xbar_mg6_wo_to_sg0_cmd_attri  [   2:   0]),
  .o0_icb_cmd_beat                (xbar_mg6_wo_to_sg0_cmd_beat   [   1:   0]),
  .o0_icb_cmd_usr                 (xbar_mg6_wo_to_sg0_cmd_usr    [   2:   0]),
  .o0_icb_rsp_ready               (xbar_mg6_wo_to_sg0_rsp_ready             ),
  .o0_icb_rsp_valid               (xbar_mg6_wo_to_sg0_rsp_valid             ),
  .o0_icb_rsp_err                 (xbar_mg6_wo_to_sg0_rsp_err               ),
  .o0_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg0_rsp_excl_ok            ),
  .o0_icb_rsp_rdata               (xbar_mg6_wo_to_sg0_rsp_rdata  [  63:   0]),
  .o0_icb_rsp_usr                 (xbar_mg6_wo_to_sg0_rsp_usr    [   2:   0]),
      .o1_icb_enable(1'b1),
      .o1_icb_cmd_valid               (xbar_mg6_wo_to_sg1_cmd_valid             ),
  .o1_icb_cmd_ready               (xbar_mg6_wo_to_sg1_cmd_ready             ),
  .o1_icb_cmd_sel                 (xbar_mg6_wo_to_sg1_cmd_sel               ),
  .o1_icb_cmd_read                (xbar_mg6_wo_to_sg1_cmd_read              ),
  .o1_icb_cmd_addr                (xbar_mg6_wo_to_sg1_cmd_addr   [  31:   0]),
  .o1_icb_cmd_wdata               (xbar_mg6_wo_to_sg1_cmd_wdata  [  63:   0]),
  .o1_icb_cmd_wmask               (xbar_mg6_wo_to_sg1_cmd_wmask  [   7:   0]),
  .o1_icb_cmd_size                (xbar_mg6_wo_to_sg1_cmd_size   [   2:   0]),
  .o1_icb_cmd_lock                (xbar_mg6_wo_to_sg1_cmd_lock              ),
  .o1_icb_cmd_excl                (xbar_mg6_wo_to_sg1_cmd_excl              ),
  .o1_icb_cmd_xlen                (xbar_mg6_wo_to_sg1_cmd_xlen   [   7:   0]),
  .o1_icb_cmd_xburst              (xbar_mg6_wo_to_sg1_cmd_xburst [   1:   0]),
  .o1_icb_cmd_modes               (xbar_mg6_wo_to_sg1_cmd_modes  [   1:   0]),
  .o1_icb_cmd_dmode               (xbar_mg6_wo_to_sg1_cmd_dmode             ),
  .o1_icb_cmd_attri               (xbar_mg6_wo_to_sg1_cmd_attri  [   2:   0]),
  .o1_icb_cmd_beat                (xbar_mg6_wo_to_sg1_cmd_beat   [   1:   0]),
  .o1_icb_cmd_usr                 (xbar_mg6_wo_to_sg1_cmd_usr    [   2:   0]),
  .o1_icb_rsp_ready               (xbar_mg6_wo_to_sg1_rsp_ready             ),
  .o1_icb_rsp_valid               (xbar_mg6_wo_to_sg1_rsp_valid             ),
  .o1_icb_rsp_err                 (xbar_mg6_wo_to_sg1_rsp_err               ),
  .o1_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg1_rsp_excl_ok            ),
  .o1_icb_rsp_rdata               (xbar_mg6_wo_to_sg1_rsp_rdata  [  63:   0]),
  .o1_icb_rsp_usr                 (xbar_mg6_wo_to_sg1_rsp_usr    [   2:   0]),
      .o2_icb_enable(1'b1),
      .o2_icb_cmd_valid               (xbar_mg6_wo_to_sg2_cmd_valid             ),
  .o2_icb_cmd_ready               (xbar_mg6_wo_to_sg2_cmd_ready             ),
  .o2_icb_cmd_sel                 (xbar_mg6_wo_to_sg2_cmd_sel               ),
  .o2_icb_cmd_read                (xbar_mg6_wo_to_sg2_cmd_read              ),
  .o2_icb_cmd_addr                (xbar_mg6_wo_to_sg2_cmd_addr   [  31:   0]),
  .o2_icb_cmd_wdata               (xbar_mg6_wo_to_sg2_cmd_wdata  [  63:   0]),
  .o2_icb_cmd_wmask               (xbar_mg6_wo_to_sg2_cmd_wmask  [   7:   0]),
  .o2_icb_cmd_size                (xbar_mg6_wo_to_sg2_cmd_size   [   2:   0]),
  .o2_icb_cmd_lock                (xbar_mg6_wo_to_sg2_cmd_lock              ),
  .o2_icb_cmd_excl                (xbar_mg6_wo_to_sg2_cmd_excl              ),
  .o2_icb_cmd_xlen                (xbar_mg6_wo_to_sg2_cmd_xlen   [   7:   0]),
  .o2_icb_cmd_xburst              (xbar_mg6_wo_to_sg2_cmd_xburst [   1:   0]),
  .o2_icb_cmd_modes               (xbar_mg6_wo_to_sg2_cmd_modes  [   1:   0]),
  .o2_icb_cmd_dmode               (xbar_mg6_wo_to_sg2_cmd_dmode             ),
  .o2_icb_cmd_attri               (xbar_mg6_wo_to_sg2_cmd_attri  [   2:   0]),
  .o2_icb_cmd_beat                (xbar_mg6_wo_to_sg2_cmd_beat   [   1:   0]),
  .o2_icb_cmd_usr                 (xbar_mg6_wo_to_sg2_cmd_usr    [   2:   0]),
  .o2_icb_rsp_ready               (xbar_mg6_wo_to_sg2_rsp_ready             ),
  .o2_icb_rsp_valid               (xbar_mg6_wo_to_sg2_rsp_valid             ),
  .o2_icb_rsp_err                 (xbar_mg6_wo_to_sg2_rsp_err               ),
  .o2_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg2_rsp_excl_ok            ),
  .o2_icb_rsp_rdata               (xbar_mg6_wo_to_sg2_rsp_rdata  [  63:   0]),
  .o2_icb_rsp_usr                 (xbar_mg6_wo_to_sg2_rsp_usr    [   2:   0]),
      .o3_icb_enable(1'b1),
      .o3_icb_cmd_valid               (xbar_mg6_wo_to_sg3_cmd_valid             ),
  .o3_icb_cmd_ready               (xbar_mg6_wo_to_sg3_cmd_ready             ),
  .o3_icb_cmd_sel                 (xbar_mg6_wo_to_sg3_cmd_sel               ),
  .o3_icb_cmd_read                (xbar_mg6_wo_to_sg3_cmd_read              ),
  .o3_icb_cmd_addr                (xbar_mg6_wo_to_sg3_cmd_addr   [  31:   0]),
  .o3_icb_cmd_wdata               (xbar_mg6_wo_to_sg3_cmd_wdata  [  63:   0]),
  .o3_icb_cmd_wmask               (xbar_mg6_wo_to_sg3_cmd_wmask  [   7:   0]),
  .o3_icb_cmd_size                (xbar_mg6_wo_to_sg3_cmd_size   [   2:   0]),
  .o3_icb_cmd_lock                (xbar_mg6_wo_to_sg3_cmd_lock              ),
  .o3_icb_cmd_excl                (xbar_mg6_wo_to_sg3_cmd_excl              ),
  .o3_icb_cmd_xlen                (xbar_mg6_wo_to_sg3_cmd_xlen   [   7:   0]),
  .o3_icb_cmd_xburst              (xbar_mg6_wo_to_sg3_cmd_xburst [   1:   0]),
  .o3_icb_cmd_modes               (xbar_mg6_wo_to_sg3_cmd_modes  [   1:   0]),
  .o3_icb_cmd_dmode               (xbar_mg6_wo_to_sg3_cmd_dmode             ),
  .o3_icb_cmd_attri               (xbar_mg6_wo_to_sg3_cmd_attri  [   2:   0]),
  .o3_icb_cmd_beat                (xbar_mg6_wo_to_sg3_cmd_beat   [   1:   0]),
  .o3_icb_cmd_usr                 (xbar_mg6_wo_to_sg3_cmd_usr    [   2:   0]),
  .o3_icb_rsp_ready               (xbar_mg6_wo_to_sg3_rsp_ready             ),
  .o3_icb_rsp_valid               (xbar_mg6_wo_to_sg3_rsp_valid             ),
  .o3_icb_rsp_err                 (xbar_mg6_wo_to_sg3_rsp_err               ),
  .o3_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg3_rsp_excl_ok            ),
  .o3_icb_rsp_rdata               (xbar_mg6_wo_to_sg3_rsp_rdata  [  63:   0]),
  .o3_icb_rsp_usr                 (xbar_mg6_wo_to_sg3_rsp_usr    [   2:   0]),
      .o4_icb_enable(1'b1),
      .o4_icb_cmd_valid               (xbar_mg6_wo_to_sg4_cmd_valid             ),
  .o4_icb_cmd_ready               (xbar_mg6_wo_to_sg4_cmd_ready             ),
  .o4_icb_cmd_sel                 (xbar_mg6_wo_to_sg4_cmd_sel               ),
  .o4_icb_cmd_read                (xbar_mg6_wo_to_sg4_cmd_read              ),
  .o4_icb_cmd_addr                (xbar_mg6_wo_to_sg4_cmd_addr   [  31:   0]),
  .o4_icb_cmd_wdata               (xbar_mg6_wo_to_sg4_cmd_wdata  [  63:   0]),
  .o4_icb_cmd_wmask               (xbar_mg6_wo_to_sg4_cmd_wmask  [   7:   0]),
  .o4_icb_cmd_size                (xbar_mg6_wo_to_sg4_cmd_size   [   2:   0]),
  .o4_icb_cmd_lock                (xbar_mg6_wo_to_sg4_cmd_lock              ),
  .o4_icb_cmd_excl                (xbar_mg6_wo_to_sg4_cmd_excl              ),
  .o4_icb_cmd_xlen                (xbar_mg6_wo_to_sg4_cmd_xlen   [   7:   0]),
  .o4_icb_cmd_xburst              (xbar_mg6_wo_to_sg4_cmd_xburst [   1:   0]),
  .o4_icb_cmd_modes               (xbar_mg6_wo_to_sg4_cmd_modes  [   1:   0]),
  .o4_icb_cmd_dmode               (xbar_mg6_wo_to_sg4_cmd_dmode             ),
  .o4_icb_cmd_attri               (xbar_mg6_wo_to_sg4_cmd_attri  [   2:   0]),
  .o4_icb_cmd_beat                (xbar_mg6_wo_to_sg4_cmd_beat   [   1:   0]),
  .o4_icb_cmd_usr                 (xbar_mg6_wo_to_sg4_cmd_usr    [   2:   0]),
  .o4_icb_rsp_ready               (xbar_mg6_wo_to_sg4_rsp_ready             ),
  .o4_icb_rsp_valid               (xbar_mg6_wo_to_sg4_rsp_valid             ),
  .o4_icb_rsp_err                 (xbar_mg6_wo_to_sg4_rsp_err               ),
  .o4_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg4_rsp_excl_ok            ),
  .o4_icb_rsp_rdata               (xbar_mg6_wo_to_sg4_rsp_rdata  [  63:   0]),
  .o4_icb_rsp_usr                 (xbar_mg6_wo_to_sg4_rsp_usr    [   2:   0]),
      .o5_icb_enable(1'b1),
      .o5_icb_cmd_valid               (xbar_mg6_wo_to_sg5_cmd_valid             ),
  .o5_icb_cmd_ready               (xbar_mg6_wo_to_sg5_cmd_ready             ),
  .o5_icb_cmd_sel                 (xbar_mg6_wo_to_sg5_cmd_sel               ),
  .o5_icb_cmd_read                (xbar_mg6_wo_to_sg5_cmd_read              ),
  .o5_icb_cmd_addr                (xbar_mg6_wo_to_sg5_cmd_addr   [  31:   0]),
  .o5_icb_cmd_wdata               (xbar_mg6_wo_to_sg5_cmd_wdata  [  63:   0]),
  .o5_icb_cmd_wmask               (xbar_mg6_wo_to_sg5_cmd_wmask  [   7:   0]),
  .o5_icb_cmd_size                (xbar_mg6_wo_to_sg5_cmd_size   [   2:   0]),
  .o5_icb_cmd_lock                (xbar_mg6_wo_to_sg5_cmd_lock              ),
  .o5_icb_cmd_excl                (xbar_mg6_wo_to_sg5_cmd_excl              ),
  .o5_icb_cmd_xlen                (xbar_mg6_wo_to_sg5_cmd_xlen   [   7:   0]),
  .o5_icb_cmd_xburst              (xbar_mg6_wo_to_sg5_cmd_xburst [   1:   0]),
  .o5_icb_cmd_modes               (xbar_mg6_wo_to_sg5_cmd_modes  [   1:   0]),
  .o5_icb_cmd_dmode               (xbar_mg6_wo_to_sg5_cmd_dmode             ),
  .o5_icb_cmd_attri               (xbar_mg6_wo_to_sg5_cmd_attri  [   2:   0]),
  .o5_icb_cmd_beat                (xbar_mg6_wo_to_sg5_cmd_beat   [   1:   0]),
  .o5_icb_cmd_usr                 (xbar_mg6_wo_to_sg5_cmd_usr    [   2:   0]),
  .o5_icb_rsp_ready               (xbar_mg6_wo_to_sg5_rsp_ready             ),
  .o5_icb_rsp_valid               (xbar_mg6_wo_to_sg5_rsp_valid             ),
  .o5_icb_rsp_err                 (xbar_mg6_wo_to_sg5_rsp_err               ),
  .o5_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg5_rsp_excl_ok            ),
  .o5_icb_rsp_rdata               (xbar_mg6_wo_to_sg5_rsp_rdata  [  63:   0]),
  .o5_icb_rsp_usr                 (xbar_mg6_wo_to_sg5_rsp_usr    [   2:   0]),
      .o6_icb_cmd_valid               (xbar_mg6_wo_to_sg6_cmd_valid             ),
  .o6_icb_cmd_ready               (xbar_mg6_wo_to_sg6_cmd_ready             ),
  .o6_icb_cmd_sel                 (xbar_mg6_wo_to_sg6_cmd_sel               ),
  .o6_icb_cmd_read                (xbar_mg6_wo_to_sg6_cmd_read              ),
  .o6_icb_cmd_addr                (xbar_mg6_wo_to_sg6_cmd_addr   [  31:   0]),
  .o6_icb_cmd_wdata               (xbar_mg6_wo_to_sg6_cmd_wdata  [  63:   0]),
  .o6_icb_cmd_wmask               (xbar_mg6_wo_to_sg6_cmd_wmask  [   7:   0]),
  .o6_icb_cmd_size                (xbar_mg6_wo_to_sg6_cmd_size   [   2:   0]),
  .o6_icb_cmd_lock                (xbar_mg6_wo_to_sg6_cmd_lock              ),
  .o6_icb_cmd_excl                (xbar_mg6_wo_to_sg6_cmd_excl              ),
  .o6_icb_cmd_xlen                (xbar_mg6_wo_to_sg6_cmd_xlen   [   7:   0]),
  .o6_icb_cmd_xburst              (xbar_mg6_wo_to_sg6_cmd_xburst [   1:   0]),
  .o6_icb_cmd_modes               (xbar_mg6_wo_to_sg6_cmd_modes  [   1:   0]),
  .o6_icb_cmd_dmode               (xbar_mg6_wo_to_sg6_cmd_dmode             ),
  .o6_icb_cmd_attri               (xbar_mg6_wo_to_sg6_cmd_attri  [   2:   0]),
  .o6_icb_cmd_beat                (xbar_mg6_wo_to_sg6_cmd_beat   [   1:   0]),
  .o6_icb_cmd_usr                 (xbar_mg6_wo_to_sg6_cmd_usr    [   2:   0]),
  .o6_icb_rsp_ready               (xbar_mg6_wo_to_sg6_rsp_ready             ),
  .o6_icb_rsp_valid               (xbar_mg6_wo_to_sg6_rsp_valid             ),
  .o6_icb_rsp_err                 (xbar_mg6_wo_to_sg6_rsp_err               ),
  .o6_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg6_rsp_excl_ok            ),
  .o6_icb_rsp_rdata               (xbar_mg6_wo_to_sg6_rsp_rdata  [  63:   0]),
  .o6_icb_rsp_usr                 (xbar_mg6_wo_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg5_ro_arbt_active;
   e603_subsys_xbar_slv5_ro_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO    (0), 
      .O_SUPPORT_RATIO    (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (128  ),
      .ARBT_FIFO_OUTS_CNT_W(8),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg5_ro_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg5_ro_arbt_active),
      .o_icb_cmd_valid                (slv_grp_5_ro_icb_cmd_valid               ),
  .o_icb_cmd_ready                (slv_grp_5_ro_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (slv_grp_5_ro_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (slv_grp_5_ro_icb_cmd_read                ),
  .o_icb_cmd_addr                 (slv_grp_5_ro_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_5_ro_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_5_ro_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_5_ro_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_5_ro_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (slv_grp_5_ro_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (slv_grp_5_ro_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_5_ro_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_5_ro_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_5_ro_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (slv_grp_5_ro_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_5_ro_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_5_ro_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_5_ro_icb_rsp_ready               ),
  .o_icb_rsp_valid                (slv_grp_5_ro_icb_rsp_valid               ),
  .o_icb_rsp_err                  (slv_grp_5_ro_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (slv_grp_5_ro_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (slv_grp_5_ro_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_5_ro_icb_rsp_usr      [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_ro_to_sg5_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_ro_to_sg5_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_ro_to_sg5_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_ro_to_sg5_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_ro_to_sg5_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_ro_to_sg5_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_ro_to_sg5_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_ro_to_sg5_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_ro_to_sg5_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_ro_to_sg5_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_ro_to_sg5_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_ro_to_sg5_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_ro_to_sg5_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_ro_to_sg5_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_ro_to_sg5_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_ro_to_sg5_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_ro_to_sg5_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_ro_to_sg5_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_ro_to_sg5_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_ro_to_sg5_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg5_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_ro_to_sg5_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_ro_to_sg5_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg1_ro_to_sg5_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg1_ro_to_sg5_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg1_ro_to_sg5_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg1_ro_to_sg5_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg1_ro_to_sg5_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg1_ro_to_sg5_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg1_ro_to_sg5_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg1_ro_to_sg5_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg1_ro_to_sg5_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg1_ro_to_sg5_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg1_ro_to_sg5_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg1_ro_to_sg5_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg1_ro_to_sg5_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg1_ro_to_sg5_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg1_ro_to_sg5_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg1_ro_to_sg5_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg1_ro_to_sg5_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg1_ro_to_sg5_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg1_ro_to_sg5_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg1_ro_to_sg5_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg5_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg1_ro_to_sg5_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg1_ro_to_sg5_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg3_ro_to_sg5_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg3_ro_to_sg5_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg3_ro_to_sg5_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg3_ro_to_sg5_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg3_ro_to_sg5_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg3_ro_to_sg5_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg3_ro_to_sg5_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg3_ro_to_sg5_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg3_ro_to_sg5_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg3_ro_to_sg5_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg3_ro_to_sg5_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg3_ro_to_sg5_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg3_ro_to_sg5_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg3_ro_to_sg5_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg3_ro_to_sg5_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg3_ro_to_sg5_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg3_ro_to_sg5_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg3_ro_to_sg5_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg3_ro_to_sg5_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg3_ro_to_sg5_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg5_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg3_ro_to_sg5_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg3_ro_to_sg5_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg4_ro_to_sg5_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg4_ro_to_sg5_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg4_ro_to_sg5_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg4_ro_to_sg5_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg4_ro_to_sg5_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg4_ro_to_sg5_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg4_ro_to_sg5_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg4_ro_to_sg5_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg4_ro_to_sg5_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg4_ro_to_sg5_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg4_ro_to_sg5_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg4_ro_to_sg5_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg4_ro_to_sg5_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg4_ro_to_sg5_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg4_ro_to_sg5_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg4_ro_to_sg5_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg4_ro_to_sg5_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg4_ro_to_sg5_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg4_ro_to_sg5_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg4_ro_to_sg5_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg5_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg4_ro_to_sg5_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg4_ro_to_sg5_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg5_ro_to_sg5_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg5_ro_to_sg5_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg5_ro_to_sg5_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg5_ro_to_sg5_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg5_ro_to_sg5_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg5_ro_to_sg5_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg5_ro_to_sg5_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg5_ro_to_sg5_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg5_ro_to_sg5_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg5_ro_to_sg5_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg5_ro_to_sg5_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg5_ro_to_sg5_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg5_ro_to_sg5_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg5_ro_to_sg5_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg5_ro_to_sg5_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg5_ro_to_sg5_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg5_ro_to_sg5_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg5_ro_to_sg5_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg5_ro_to_sg5_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg5_ro_to_sg5_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg5_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg5_ro_to_sg5_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg5_ro_to_sg5_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg6_ro_to_sg5_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg6_ro_to_sg5_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg6_ro_to_sg5_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg6_ro_to_sg5_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg6_ro_to_sg5_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg6_ro_to_sg5_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg6_ro_to_sg5_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg6_ro_to_sg5_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg6_ro_to_sg5_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg6_ro_to_sg5_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg6_ro_to_sg5_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg6_ro_to_sg5_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg6_ro_to_sg5_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg6_ro_to_sg5_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg6_ro_to_sg5_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg6_ro_to_sg5_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg6_ro_to_sg5_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg6_ro_to_sg5_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg6_ro_to_sg5_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg6_ro_to_sg5_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg6_ro_to_sg5_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg6_ro_to_sg5_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg6_ro_to_sg5_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg5_wo_arbt_active;
   e603_subsys_xbar_slv5_wo_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO    (0), 
      .O_SUPPORT_RATIO    (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (128  ),
      .ARBT_FIFO_OUTS_CNT_W(8),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg5_wo_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg5_wo_arbt_active),
      .o_icb_cmd_valid                (slv_grp_5_wo_icb_cmd_valid               ),
  .o_icb_cmd_ready                (slv_grp_5_wo_icb_cmd_ready               ),
  .o_icb_cmd_sel                  (slv_grp_5_wo_icb_cmd_sel                 ),
  .o_icb_cmd_read                 (slv_grp_5_wo_icb_cmd_read                ),
  .o_icb_cmd_addr                 (slv_grp_5_wo_icb_cmd_addr     [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_5_wo_icb_cmd_wdata    [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_5_wo_icb_cmd_wmask    [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_5_wo_icb_cmd_size     [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_5_wo_icb_cmd_lock                ),
  .o_icb_cmd_excl                 (slv_grp_5_wo_icb_cmd_excl                ),
  .o_icb_cmd_xlen                 (slv_grp_5_wo_icb_cmd_xlen     [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_5_wo_icb_cmd_xburst   [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_5_wo_icb_cmd_modes    [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_5_wo_icb_cmd_dmode               ),
  .o_icb_cmd_attri                (slv_grp_5_wo_icb_cmd_attri    [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_5_wo_icb_cmd_beat     [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_5_wo_icb_cmd_usr      [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_5_wo_icb_rsp_ready               ),
  .o_icb_rsp_valid                (slv_grp_5_wo_icb_rsp_valid               ),
  .o_icb_rsp_err                  (slv_grp_5_wo_icb_rsp_err                 ),
  .o_icb_rsp_excl_ok              (slv_grp_5_wo_icb_rsp_excl_ok             ),
  .o_icb_rsp_rdata                (slv_grp_5_wo_icb_rsp_rdata    [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_5_wo_icb_rsp_usr      [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_wo_to_sg5_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_wo_to_sg5_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_wo_to_sg5_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_wo_to_sg5_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_wo_to_sg5_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_wo_to_sg5_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_wo_to_sg5_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_wo_to_sg5_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_wo_to_sg5_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_wo_to_sg5_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_wo_to_sg5_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_wo_to_sg5_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_wo_to_sg5_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_wo_to_sg5_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_wo_to_sg5_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_wo_to_sg5_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_wo_to_sg5_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_wo_to_sg5_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_wo_to_sg5_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_wo_to_sg5_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg5_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_wo_to_sg5_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_wo_to_sg5_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg2_wo_to_sg5_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg2_wo_to_sg5_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg2_wo_to_sg5_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg2_wo_to_sg5_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg2_wo_to_sg5_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg2_wo_to_sg5_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg2_wo_to_sg5_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg2_wo_to_sg5_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg2_wo_to_sg5_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg2_wo_to_sg5_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg2_wo_to_sg5_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg2_wo_to_sg5_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg2_wo_to_sg5_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg2_wo_to_sg5_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg2_wo_to_sg5_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg2_wo_to_sg5_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg2_wo_to_sg5_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg2_wo_to_sg5_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg2_wo_to_sg5_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg2_wo_to_sg5_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg5_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg2_wo_to_sg5_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg2_wo_to_sg5_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg3_wo_to_sg5_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg3_wo_to_sg5_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg3_wo_to_sg5_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg3_wo_to_sg5_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg3_wo_to_sg5_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg3_wo_to_sg5_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg3_wo_to_sg5_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg3_wo_to_sg5_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg3_wo_to_sg5_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg3_wo_to_sg5_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg3_wo_to_sg5_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg3_wo_to_sg5_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg3_wo_to_sg5_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg3_wo_to_sg5_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg3_wo_to_sg5_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg3_wo_to_sg5_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg3_wo_to_sg5_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg3_wo_to_sg5_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg3_wo_to_sg5_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg3_wo_to_sg5_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg5_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg3_wo_to_sg5_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg3_wo_to_sg5_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg4_wo_to_sg5_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg4_wo_to_sg5_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg4_wo_to_sg5_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg4_wo_to_sg5_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg4_wo_to_sg5_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg4_wo_to_sg5_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg4_wo_to_sg5_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg4_wo_to_sg5_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg4_wo_to_sg5_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg4_wo_to_sg5_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg4_wo_to_sg5_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg4_wo_to_sg5_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg4_wo_to_sg5_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg4_wo_to_sg5_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg4_wo_to_sg5_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg4_wo_to_sg5_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg4_wo_to_sg5_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg4_wo_to_sg5_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg4_wo_to_sg5_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg4_wo_to_sg5_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg5_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg4_wo_to_sg5_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg4_wo_to_sg5_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg5_wo_to_sg5_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg5_wo_to_sg5_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg5_wo_to_sg5_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg5_wo_to_sg5_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg5_wo_to_sg5_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg5_wo_to_sg5_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg5_wo_to_sg5_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg5_wo_to_sg5_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg5_wo_to_sg5_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg5_wo_to_sg5_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg5_wo_to_sg5_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg5_wo_to_sg5_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg5_wo_to_sg5_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg5_wo_to_sg5_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg5_wo_to_sg5_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg5_wo_to_sg5_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg5_wo_to_sg5_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg5_wo_to_sg5_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg5_wo_to_sg5_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg5_wo_to_sg5_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg5_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg5_wo_to_sg5_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg5_wo_to_sg5_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg6_wo_to_sg5_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg6_wo_to_sg5_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg6_wo_to_sg5_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg6_wo_to_sg5_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg6_wo_to_sg5_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg6_wo_to_sg5_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg6_wo_to_sg5_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg6_wo_to_sg5_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg6_wo_to_sg5_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg6_wo_to_sg5_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg6_wo_to_sg5_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg6_wo_to_sg5_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg6_wo_to_sg5_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg6_wo_to_sg5_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg6_wo_to_sg5_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg6_wo_to_sg5_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg6_wo_to_sg5_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg6_wo_to_sg5_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg6_wo_to_sg5_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg6_wo_to_sg5_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg6_wo_to_sg5_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg6_wo_to_sg5_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg6_wo_to_sg5_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg0_rw_arbt_active;
   e603_subsys_xbar_slv0_rw_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (16  ),
      .ARBT_FIFO_OUTS_CNT_W(5),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg0_rw_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg0_rw_arbt_active),
      .o_icb_cmd_valid                (slv_grp_0_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (slv_grp_0_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (slv_grp_0_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (slv_grp_0_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (slv_grp_0_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_0_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_0_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_0_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_0_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (slv_grp_0_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (slv_grp_0_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_0_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_0_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_0_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (slv_grp_0_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_0_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_0_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_0_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (slv_grp_0_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (slv_grp_0_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (slv_grp_0_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (slv_grp_0_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_0_icb_rsp_usr         [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_ro_to_sg0_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_ro_to_sg0_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_ro_to_sg0_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_ro_to_sg0_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_ro_to_sg0_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_ro_to_sg0_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_ro_to_sg0_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_ro_to_sg0_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_ro_to_sg0_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_ro_to_sg0_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_ro_to_sg0_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_ro_to_sg0_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_ro_to_sg0_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_ro_to_sg0_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_ro_to_sg0_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_ro_to_sg0_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_ro_to_sg0_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_ro_to_sg0_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_ro_to_sg0_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_ro_to_sg0_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg0_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_ro_to_sg0_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_ro_to_sg0_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg0_wo_to_sg0_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg0_wo_to_sg0_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg0_wo_to_sg0_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg0_wo_to_sg0_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg0_wo_to_sg0_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg0_wo_to_sg0_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg0_wo_to_sg0_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg0_wo_to_sg0_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg0_wo_to_sg0_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg0_wo_to_sg0_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg0_wo_to_sg0_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg0_wo_to_sg0_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg0_wo_to_sg0_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg0_wo_to_sg0_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg0_wo_to_sg0_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg0_wo_to_sg0_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg0_wo_to_sg0_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg0_wo_to_sg0_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg0_wo_to_sg0_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg0_wo_to_sg0_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg0_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg0_wo_to_sg0_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg0_wo_to_sg0_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg1_ro_to_sg0_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg1_ro_to_sg0_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg1_ro_to_sg0_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg1_ro_to_sg0_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg1_ro_to_sg0_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg1_ro_to_sg0_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg1_ro_to_sg0_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg1_ro_to_sg0_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg1_ro_to_sg0_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg1_ro_to_sg0_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg1_ro_to_sg0_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg1_ro_to_sg0_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg1_ro_to_sg0_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg1_ro_to_sg0_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg1_ro_to_sg0_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg1_ro_to_sg0_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg1_ro_to_sg0_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg1_ro_to_sg0_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg1_ro_to_sg0_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg1_ro_to_sg0_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg0_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg1_ro_to_sg0_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg1_ro_to_sg0_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg2_wo_to_sg0_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg2_wo_to_sg0_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg2_wo_to_sg0_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg2_wo_to_sg0_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg2_wo_to_sg0_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg2_wo_to_sg0_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg2_wo_to_sg0_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg2_wo_to_sg0_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg2_wo_to_sg0_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg2_wo_to_sg0_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg2_wo_to_sg0_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg2_wo_to_sg0_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg2_wo_to_sg0_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg2_wo_to_sg0_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg2_wo_to_sg0_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg2_wo_to_sg0_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg2_wo_to_sg0_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg2_wo_to_sg0_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg2_wo_to_sg0_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg2_wo_to_sg0_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg0_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg2_wo_to_sg0_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg2_wo_to_sg0_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg3_ro_to_sg0_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg3_ro_to_sg0_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg3_ro_to_sg0_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg3_ro_to_sg0_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg3_ro_to_sg0_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg3_ro_to_sg0_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg3_ro_to_sg0_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg3_ro_to_sg0_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg3_ro_to_sg0_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg3_ro_to_sg0_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg3_ro_to_sg0_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg3_ro_to_sg0_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg3_ro_to_sg0_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg3_ro_to_sg0_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg3_ro_to_sg0_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg3_ro_to_sg0_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg3_ro_to_sg0_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg3_ro_to_sg0_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg3_ro_to_sg0_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg3_ro_to_sg0_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg0_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg3_ro_to_sg0_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg3_ro_to_sg0_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg3_wo_to_sg0_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg3_wo_to_sg0_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg3_wo_to_sg0_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg3_wo_to_sg0_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg3_wo_to_sg0_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg3_wo_to_sg0_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg3_wo_to_sg0_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg3_wo_to_sg0_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg3_wo_to_sg0_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg3_wo_to_sg0_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg3_wo_to_sg0_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg3_wo_to_sg0_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg3_wo_to_sg0_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg3_wo_to_sg0_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg3_wo_to_sg0_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg3_wo_to_sg0_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg3_wo_to_sg0_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg3_wo_to_sg0_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg3_wo_to_sg0_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg3_wo_to_sg0_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg0_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg3_wo_to_sg0_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg3_wo_to_sg0_rsp_usr    [   2:   0]),
      .i6_icb_cmd_valid               (xbar_mg4_ro_to_sg0_cmd_valid             ),
  .i6_icb_cmd_ready               (xbar_mg4_ro_to_sg0_cmd_ready             ),
  .i6_icb_cmd_sel                 (xbar_mg4_ro_to_sg0_cmd_sel               ),
  .i6_icb_cmd_read                (xbar_mg4_ro_to_sg0_cmd_read              ),
  .i6_icb_cmd_addr                (xbar_mg4_ro_to_sg0_cmd_addr   [  31:   0]),
  .i6_icb_cmd_wdata               (xbar_mg4_ro_to_sg0_cmd_wdata  [  63:   0]),
  .i6_icb_cmd_wmask               (xbar_mg4_ro_to_sg0_cmd_wmask  [   7:   0]),
  .i6_icb_cmd_size                (xbar_mg4_ro_to_sg0_cmd_size   [   2:   0]),
  .i6_icb_cmd_lock                (xbar_mg4_ro_to_sg0_cmd_lock              ),
  .i6_icb_cmd_excl                (xbar_mg4_ro_to_sg0_cmd_excl              ),
  .i6_icb_cmd_xlen                (xbar_mg4_ro_to_sg0_cmd_xlen   [   7:   0]),
  .i6_icb_cmd_xburst              (xbar_mg4_ro_to_sg0_cmd_xburst [   1:   0]),
  .i6_icb_cmd_modes               (xbar_mg4_ro_to_sg0_cmd_modes  [   1:   0]),
  .i6_icb_cmd_dmode               (xbar_mg4_ro_to_sg0_cmd_dmode             ),
  .i6_icb_cmd_attri               (xbar_mg4_ro_to_sg0_cmd_attri  [   2:   0]),
  .i6_icb_cmd_beat                (xbar_mg4_ro_to_sg0_cmd_beat   [   1:   0]),
  .i6_icb_cmd_usr                 (xbar_mg4_ro_to_sg0_cmd_usr    [   2:   0]),
  .i6_icb_rsp_ready               (xbar_mg4_ro_to_sg0_rsp_ready             ),
  .i6_icb_rsp_valid               (xbar_mg4_ro_to_sg0_rsp_valid             ),
  .i6_icb_rsp_err                 (xbar_mg4_ro_to_sg0_rsp_err               ),
  .i6_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg0_rsp_excl_ok            ),
  .i6_icb_rsp_rdata               (xbar_mg4_ro_to_sg0_rsp_rdata  [  63:   0]),
  .i6_icb_rsp_usr                 (xbar_mg4_ro_to_sg0_rsp_usr    [   2:   0]),
      .i7_icb_cmd_valid               (xbar_mg4_wo_to_sg0_cmd_valid             ),
  .i7_icb_cmd_ready               (xbar_mg4_wo_to_sg0_cmd_ready             ),
  .i7_icb_cmd_sel                 (xbar_mg4_wo_to_sg0_cmd_sel               ),
  .i7_icb_cmd_read                (xbar_mg4_wo_to_sg0_cmd_read              ),
  .i7_icb_cmd_addr                (xbar_mg4_wo_to_sg0_cmd_addr   [  31:   0]),
  .i7_icb_cmd_wdata               (xbar_mg4_wo_to_sg0_cmd_wdata  [  63:   0]),
  .i7_icb_cmd_wmask               (xbar_mg4_wo_to_sg0_cmd_wmask  [   7:   0]),
  .i7_icb_cmd_size                (xbar_mg4_wo_to_sg0_cmd_size   [   2:   0]),
  .i7_icb_cmd_lock                (xbar_mg4_wo_to_sg0_cmd_lock              ),
  .i7_icb_cmd_excl                (xbar_mg4_wo_to_sg0_cmd_excl              ),
  .i7_icb_cmd_xlen                (xbar_mg4_wo_to_sg0_cmd_xlen   [   7:   0]),
  .i7_icb_cmd_xburst              (xbar_mg4_wo_to_sg0_cmd_xburst [   1:   0]),
  .i7_icb_cmd_modes               (xbar_mg4_wo_to_sg0_cmd_modes  [   1:   0]),
  .i7_icb_cmd_dmode               (xbar_mg4_wo_to_sg0_cmd_dmode             ),
  .i7_icb_cmd_attri               (xbar_mg4_wo_to_sg0_cmd_attri  [   2:   0]),
  .i7_icb_cmd_beat                (xbar_mg4_wo_to_sg0_cmd_beat   [   1:   0]),
  .i7_icb_cmd_usr                 (xbar_mg4_wo_to_sg0_cmd_usr    [   2:   0]),
  .i7_icb_rsp_ready               (xbar_mg4_wo_to_sg0_rsp_ready             ),
  .i7_icb_rsp_valid               (xbar_mg4_wo_to_sg0_rsp_valid             ),
  .i7_icb_rsp_err                 (xbar_mg4_wo_to_sg0_rsp_err               ),
  .i7_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg0_rsp_excl_ok            ),
  .i7_icb_rsp_rdata               (xbar_mg4_wo_to_sg0_rsp_rdata  [  63:   0]),
  .i7_icb_rsp_usr                 (xbar_mg4_wo_to_sg0_rsp_usr    [   2:   0]),
      .i8_icb_cmd_valid               (xbar_mg5_ro_to_sg0_cmd_valid             ),
  .i8_icb_cmd_ready               (xbar_mg5_ro_to_sg0_cmd_ready             ),
  .i8_icb_cmd_sel                 (xbar_mg5_ro_to_sg0_cmd_sel               ),
  .i8_icb_cmd_read                (xbar_mg5_ro_to_sg0_cmd_read              ),
  .i8_icb_cmd_addr                (xbar_mg5_ro_to_sg0_cmd_addr   [  31:   0]),
  .i8_icb_cmd_wdata               (xbar_mg5_ro_to_sg0_cmd_wdata  [  63:   0]),
  .i8_icb_cmd_wmask               (xbar_mg5_ro_to_sg0_cmd_wmask  [   7:   0]),
  .i8_icb_cmd_size                (xbar_mg5_ro_to_sg0_cmd_size   [   2:   0]),
  .i8_icb_cmd_lock                (xbar_mg5_ro_to_sg0_cmd_lock              ),
  .i8_icb_cmd_excl                (xbar_mg5_ro_to_sg0_cmd_excl              ),
  .i8_icb_cmd_xlen                (xbar_mg5_ro_to_sg0_cmd_xlen   [   7:   0]),
  .i8_icb_cmd_xburst              (xbar_mg5_ro_to_sg0_cmd_xburst [   1:   0]),
  .i8_icb_cmd_modes               (xbar_mg5_ro_to_sg0_cmd_modes  [   1:   0]),
  .i8_icb_cmd_dmode               (xbar_mg5_ro_to_sg0_cmd_dmode             ),
  .i8_icb_cmd_attri               (xbar_mg5_ro_to_sg0_cmd_attri  [   2:   0]),
  .i8_icb_cmd_beat                (xbar_mg5_ro_to_sg0_cmd_beat   [   1:   0]),
  .i8_icb_cmd_usr                 (xbar_mg5_ro_to_sg0_cmd_usr    [   2:   0]),
  .i8_icb_rsp_ready               (xbar_mg5_ro_to_sg0_rsp_ready             ),
  .i8_icb_rsp_valid               (xbar_mg5_ro_to_sg0_rsp_valid             ),
  .i8_icb_rsp_err                 (xbar_mg5_ro_to_sg0_rsp_err               ),
  .i8_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg0_rsp_excl_ok            ),
  .i8_icb_rsp_rdata               (xbar_mg5_ro_to_sg0_rsp_rdata  [  63:   0]),
  .i8_icb_rsp_usr                 (xbar_mg5_ro_to_sg0_rsp_usr    [   2:   0]),
      .i9_icb_cmd_valid               (xbar_mg5_wo_to_sg0_cmd_valid             ),
  .i9_icb_cmd_ready               (xbar_mg5_wo_to_sg0_cmd_ready             ),
  .i9_icb_cmd_sel                 (xbar_mg5_wo_to_sg0_cmd_sel               ),
  .i9_icb_cmd_read                (xbar_mg5_wo_to_sg0_cmd_read              ),
  .i9_icb_cmd_addr                (xbar_mg5_wo_to_sg0_cmd_addr   [  31:   0]),
  .i9_icb_cmd_wdata               (xbar_mg5_wo_to_sg0_cmd_wdata  [  63:   0]),
  .i9_icb_cmd_wmask               (xbar_mg5_wo_to_sg0_cmd_wmask  [   7:   0]),
  .i9_icb_cmd_size                (xbar_mg5_wo_to_sg0_cmd_size   [   2:   0]),
  .i9_icb_cmd_lock                (xbar_mg5_wo_to_sg0_cmd_lock              ),
  .i9_icb_cmd_excl                (xbar_mg5_wo_to_sg0_cmd_excl              ),
  .i9_icb_cmd_xlen                (xbar_mg5_wo_to_sg0_cmd_xlen   [   7:   0]),
  .i9_icb_cmd_xburst              (xbar_mg5_wo_to_sg0_cmd_xburst [   1:   0]),
  .i9_icb_cmd_modes               (xbar_mg5_wo_to_sg0_cmd_modes  [   1:   0]),
  .i9_icb_cmd_dmode               (xbar_mg5_wo_to_sg0_cmd_dmode             ),
  .i9_icb_cmd_attri               (xbar_mg5_wo_to_sg0_cmd_attri  [   2:   0]),
  .i9_icb_cmd_beat                (xbar_mg5_wo_to_sg0_cmd_beat   [   1:   0]),
  .i9_icb_cmd_usr                 (xbar_mg5_wo_to_sg0_cmd_usr    [   2:   0]),
  .i9_icb_rsp_ready               (xbar_mg5_wo_to_sg0_rsp_ready             ),
  .i9_icb_rsp_valid               (xbar_mg5_wo_to_sg0_rsp_valid             ),
  .i9_icb_rsp_err                 (xbar_mg5_wo_to_sg0_rsp_err               ),
  .i9_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg0_rsp_excl_ok            ),
  .i9_icb_rsp_rdata               (xbar_mg5_wo_to_sg0_rsp_rdata  [  63:   0]),
  .i9_icb_rsp_usr                 (xbar_mg5_wo_to_sg0_rsp_usr    [   2:   0]),
      .i10_icb_cmd_valid              (xbar_mg6_ro_to_sg0_cmd_valid             ),
  .i10_icb_cmd_ready              (xbar_mg6_ro_to_sg0_cmd_ready             ),
  .i10_icb_cmd_sel                (xbar_mg6_ro_to_sg0_cmd_sel               ),
  .i10_icb_cmd_read               (xbar_mg6_ro_to_sg0_cmd_read              ),
  .i10_icb_cmd_addr               (xbar_mg6_ro_to_sg0_cmd_addr   [  31:   0]),
  .i10_icb_cmd_wdata              (xbar_mg6_ro_to_sg0_cmd_wdata  [  63:   0]),
  .i10_icb_cmd_wmask              (xbar_mg6_ro_to_sg0_cmd_wmask  [   7:   0]),
  .i10_icb_cmd_size               (xbar_mg6_ro_to_sg0_cmd_size   [   2:   0]),
  .i10_icb_cmd_lock               (xbar_mg6_ro_to_sg0_cmd_lock              ),
  .i10_icb_cmd_excl               (xbar_mg6_ro_to_sg0_cmd_excl              ),
  .i10_icb_cmd_xlen               (xbar_mg6_ro_to_sg0_cmd_xlen   [   7:   0]),
  .i10_icb_cmd_xburst             (xbar_mg6_ro_to_sg0_cmd_xburst [   1:   0]),
  .i10_icb_cmd_modes              (xbar_mg6_ro_to_sg0_cmd_modes  [   1:   0]),
  .i10_icb_cmd_dmode              (xbar_mg6_ro_to_sg0_cmd_dmode             ),
  .i10_icb_cmd_attri              (xbar_mg6_ro_to_sg0_cmd_attri  [   2:   0]),
  .i10_icb_cmd_beat               (xbar_mg6_ro_to_sg0_cmd_beat   [   1:   0]),
  .i10_icb_cmd_usr                (xbar_mg6_ro_to_sg0_cmd_usr    [   2:   0]),
  .i10_icb_rsp_ready              (xbar_mg6_ro_to_sg0_rsp_ready             ),
  .i10_icb_rsp_valid              (xbar_mg6_ro_to_sg0_rsp_valid             ),
  .i10_icb_rsp_err                (xbar_mg6_ro_to_sg0_rsp_err               ),
  .i10_icb_rsp_excl_ok            (xbar_mg6_ro_to_sg0_rsp_excl_ok            ),
  .i10_icb_rsp_rdata              (xbar_mg6_ro_to_sg0_rsp_rdata  [  63:   0]),
  .i10_icb_rsp_usr                (xbar_mg6_ro_to_sg0_rsp_usr    [   2:   0]),
      .i11_icb_cmd_valid              (xbar_mg6_wo_to_sg0_cmd_valid             ),
  .i11_icb_cmd_ready              (xbar_mg6_wo_to_sg0_cmd_ready             ),
  .i11_icb_cmd_sel                (xbar_mg6_wo_to_sg0_cmd_sel               ),
  .i11_icb_cmd_read               (xbar_mg6_wo_to_sg0_cmd_read              ),
  .i11_icb_cmd_addr               (xbar_mg6_wo_to_sg0_cmd_addr   [  31:   0]),
  .i11_icb_cmd_wdata              (xbar_mg6_wo_to_sg0_cmd_wdata  [  63:   0]),
  .i11_icb_cmd_wmask              (xbar_mg6_wo_to_sg0_cmd_wmask  [   7:   0]),
  .i11_icb_cmd_size               (xbar_mg6_wo_to_sg0_cmd_size   [   2:   0]),
  .i11_icb_cmd_lock               (xbar_mg6_wo_to_sg0_cmd_lock              ),
  .i11_icb_cmd_excl               (xbar_mg6_wo_to_sg0_cmd_excl              ),
  .i11_icb_cmd_xlen               (xbar_mg6_wo_to_sg0_cmd_xlen   [   7:   0]),
  .i11_icb_cmd_xburst             (xbar_mg6_wo_to_sg0_cmd_xburst [   1:   0]),
  .i11_icb_cmd_modes              (xbar_mg6_wo_to_sg0_cmd_modes  [   1:   0]),
  .i11_icb_cmd_dmode              (xbar_mg6_wo_to_sg0_cmd_dmode             ),
  .i11_icb_cmd_attri              (xbar_mg6_wo_to_sg0_cmd_attri  [   2:   0]),
  .i11_icb_cmd_beat               (xbar_mg6_wo_to_sg0_cmd_beat   [   1:   0]),
  .i11_icb_cmd_usr                (xbar_mg6_wo_to_sg0_cmd_usr    [   2:   0]),
  .i11_icb_rsp_ready              (xbar_mg6_wo_to_sg0_rsp_ready             ),
  .i11_icb_rsp_valid              (xbar_mg6_wo_to_sg0_rsp_valid             ),
  .i11_icb_rsp_err                (xbar_mg6_wo_to_sg0_rsp_err               ),
  .i11_icb_rsp_excl_ok            (xbar_mg6_wo_to_sg0_rsp_excl_ok            ),
  .i11_icb_rsp_rdata              (xbar_mg6_wo_to_sg0_rsp_rdata  [  63:   0]),
  .i11_icb_rsp_usr                (xbar_mg6_wo_to_sg0_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg1_rw_arbt_active;
   e603_subsys_xbar_slv1_rw_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (16  ),
      .ARBT_FIFO_OUTS_CNT_W(5),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg1_rw_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg1_rw_arbt_active),
      .o_icb_cmd_valid                (slv_grp_1_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (slv_grp_1_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (slv_grp_1_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (slv_grp_1_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (slv_grp_1_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_1_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_1_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_1_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_1_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (slv_grp_1_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (slv_grp_1_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_1_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_1_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_1_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (slv_grp_1_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_1_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_1_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_1_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (slv_grp_1_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (slv_grp_1_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (slv_grp_1_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (slv_grp_1_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_1_icb_rsp_usr         [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_ro_to_sg1_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_ro_to_sg1_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_ro_to_sg1_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_ro_to_sg1_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_ro_to_sg1_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_ro_to_sg1_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_ro_to_sg1_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_ro_to_sg1_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_ro_to_sg1_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_ro_to_sg1_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_ro_to_sg1_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_ro_to_sg1_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_ro_to_sg1_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_ro_to_sg1_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_ro_to_sg1_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_ro_to_sg1_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_ro_to_sg1_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_ro_to_sg1_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_ro_to_sg1_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_ro_to_sg1_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg1_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_ro_to_sg1_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_ro_to_sg1_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg0_wo_to_sg1_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg0_wo_to_sg1_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg0_wo_to_sg1_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg0_wo_to_sg1_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg0_wo_to_sg1_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg0_wo_to_sg1_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg0_wo_to_sg1_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg0_wo_to_sg1_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg0_wo_to_sg1_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg0_wo_to_sg1_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg0_wo_to_sg1_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg0_wo_to_sg1_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg0_wo_to_sg1_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg0_wo_to_sg1_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg0_wo_to_sg1_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg0_wo_to_sg1_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg0_wo_to_sg1_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg0_wo_to_sg1_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg0_wo_to_sg1_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg0_wo_to_sg1_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg1_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg0_wo_to_sg1_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg0_wo_to_sg1_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg1_ro_to_sg1_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg1_ro_to_sg1_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg1_ro_to_sg1_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg1_ro_to_sg1_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg1_ro_to_sg1_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg1_ro_to_sg1_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg1_ro_to_sg1_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg1_ro_to_sg1_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg1_ro_to_sg1_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg1_ro_to_sg1_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg1_ro_to_sg1_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg1_ro_to_sg1_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg1_ro_to_sg1_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg1_ro_to_sg1_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg1_ro_to_sg1_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg1_ro_to_sg1_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg1_ro_to_sg1_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg1_ro_to_sg1_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg1_ro_to_sg1_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg1_ro_to_sg1_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg1_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg1_ro_to_sg1_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg1_ro_to_sg1_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg2_wo_to_sg1_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg2_wo_to_sg1_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg2_wo_to_sg1_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg2_wo_to_sg1_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg2_wo_to_sg1_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg2_wo_to_sg1_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg2_wo_to_sg1_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg2_wo_to_sg1_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg2_wo_to_sg1_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg2_wo_to_sg1_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg2_wo_to_sg1_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg2_wo_to_sg1_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg2_wo_to_sg1_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg2_wo_to_sg1_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg2_wo_to_sg1_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg2_wo_to_sg1_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg2_wo_to_sg1_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg2_wo_to_sg1_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg2_wo_to_sg1_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg2_wo_to_sg1_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg1_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg2_wo_to_sg1_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg2_wo_to_sg1_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg3_ro_to_sg1_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg3_ro_to_sg1_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg3_ro_to_sg1_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg3_ro_to_sg1_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg3_ro_to_sg1_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg3_ro_to_sg1_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg3_ro_to_sg1_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg3_ro_to_sg1_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg3_ro_to_sg1_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg3_ro_to_sg1_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg3_ro_to_sg1_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg3_ro_to_sg1_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg3_ro_to_sg1_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg3_ro_to_sg1_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg3_ro_to_sg1_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg3_ro_to_sg1_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg3_ro_to_sg1_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg3_ro_to_sg1_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg3_ro_to_sg1_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg3_ro_to_sg1_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg1_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg3_ro_to_sg1_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg3_ro_to_sg1_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg3_wo_to_sg1_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg3_wo_to_sg1_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg3_wo_to_sg1_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg3_wo_to_sg1_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg3_wo_to_sg1_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg3_wo_to_sg1_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg3_wo_to_sg1_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg3_wo_to_sg1_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg3_wo_to_sg1_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg3_wo_to_sg1_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg3_wo_to_sg1_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg3_wo_to_sg1_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg3_wo_to_sg1_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg3_wo_to_sg1_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg3_wo_to_sg1_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg3_wo_to_sg1_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg3_wo_to_sg1_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg3_wo_to_sg1_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg3_wo_to_sg1_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg3_wo_to_sg1_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg1_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg3_wo_to_sg1_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg3_wo_to_sg1_rsp_usr    [   2:   0]),
      .i6_icb_cmd_valid               (xbar_mg4_ro_to_sg1_cmd_valid             ),
  .i6_icb_cmd_ready               (xbar_mg4_ro_to_sg1_cmd_ready             ),
  .i6_icb_cmd_sel                 (xbar_mg4_ro_to_sg1_cmd_sel               ),
  .i6_icb_cmd_read                (xbar_mg4_ro_to_sg1_cmd_read              ),
  .i6_icb_cmd_addr                (xbar_mg4_ro_to_sg1_cmd_addr   [  31:   0]),
  .i6_icb_cmd_wdata               (xbar_mg4_ro_to_sg1_cmd_wdata  [  63:   0]),
  .i6_icb_cmd_wmask               (xbar_mg4_ro_to_sg1_cmd_wmask  [   7:   0]),
  .i6_icb_cmd_size                (xbar_mg4_ro_to_sg1_cmd_size   [   2:   0]),
  .i6_icb_cmd_lock                (xbar_mg4_ro_to_sg1_cmd_lock              ),
  .i6_icb_cmd_excl                (xbar_mg4_ro_to_sg1_cmd_excl              ),
  .i6_icb_cmd_xlen                (xbar_mg4_ro_to_sg1_cmd_xlen   [   7:   0]),
  .i6_icb_cmd_xburst              (xbar_mg4_ro_to_sg1_cmd_xburst [   1:   0]),
  .i6_icb_cmd_modes               (xbar_mg4_ro_to_sg1_cmd_modes  [   1:   0]),
  .i6_icb_cmd_dmode               (xbar_mg4_ro_to_sg1_cmd_dmode             ),
  .i6_icb_cmd_attri               (xbar_mg4_ro_to_sg1_cmd_attri  [   2:   0]),
  .i6_icb_cmd_beat                (xbar_mg4_ro_to_sg1_cmd_beat   [   1:   0]),
  .i6_icb_cmd_usr                 (xbar_mg4_ro_to_sg1_cmd_usr    [   2:   0]),
  .i6_icb_rsp_ready               (xbar_mg4_ro_to_sg1_rsp_ready             ),
  .i6_icb_rsp_valid               (xbar_mg4_ro_to_sg1_rsp_valid             ),
  .i6_icb_rsp_err                 (xbar_mg4_ro_to_sg1_rsp_err               ),
  .i6_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg1_rsp_excl_ok            ),
  .i6_icb_rsp_rdata               (xbar_mg4_ro_to_sg1_rsp_rdata  [  63:   0]),
  .i6_icb_rsp_usr                 (xbar_mg4_ro_to_sg1_rsp_usr    [   2:   0]),
      .i7_icb_cmd_valid               (xbar_mg4_wo_to_sg1_cmd_valid             ),
  .i7_icb_cmd_ready               (xbar_mg4_wo_to_sg1_cmd_ready             ),
  .i7_icb_cmd_sel                 (xbar_mg4_wo_to_sg1_cmd_sel               ),
  .i7_icb_cmd_read                (xbar_mg4_wo_to_sg1_cmd_read              ),
  .i7_icb_cmd_addr                (xbar_mg4_wo_to_sg1_cmd_addr   [  31:   0]),
  .i7_icb_cmd_wdata               (xbar_mg4_wo_to_sg1_cmd_wdata  [  63:   0]),
  .i7_icb_cmd_wmask               (xbar_mg4_wo_to_sg1_cmd_wmask  [   7:   0]),
  .i7_icb_cmd_size                (xbar_mg4_wo_to_sg1_cmd_size   [   2:   0]),
  .i7_icb_cmd_lock                (xbar_mg4_wo_to_sg1_cmd_lock              ),
  .i7_icb_cmd_excl                (xbar_mg4_wo_to_sg1_cmd_excl              ),
  .i7_icb_cmd_xlen                (xbar_mg4_wo_to_sg1_cmd_xlen   [   7:   0]),
  .i7_icb_cmd_xburst              (xbar_mg4_wo_to_sg1_cmd_xburst [   1:   0]),
  .i7_icb_cmd_modes               (xbar_mg4_wo_to_sg1_cmd_modes  [   1:   0]),
  .i7_icb_cmd_dmode               (xbar_mg4_wo_to_sg1_cmd_dmode             ),
  .i7_icb_cmd_attri               (xbar_mg4_wo_to_sg1_cmd_attri  [   2:   0]),
  .i7_icb_cmd_beat                (xbar_mg4_wo_to_sg1_cmd_beat   [   1:   0]),
  .i7_icb_cmd_usr                 (xbar_mg4_wo_to_sg1_cmd_usr    [   2:   0]),
  .i7_icb_rsp_ready               (xbar_mg4_wo_to_sg1_rsp_ready             ),
  .i7_icb_rsp_valid               (xbar_mg4_wo_to_sg1_rsp_valid             ),
  .i7_icb_rsp_err                 (xbar_mg4_wo_to_sg1_rsp_err               ),
  .i7_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg1_rsp_excl_ok            ),
  .i7_icb_rsp_rdata               (xbar_mg4_wo_to_sg1_rsp_rdata  [  63:   0]),
  .i7_icb_rsp_usr                 (xbar_mg4_wo_to_sg1_rsp_usr    [   2:   0]),
      .i8_icb_cmd_valid               (xbar_mg5_ro_to_sg1_cmd_valid             ),
  .i8_icb_cmd_ready               (xbar_mg5_ro_to_sg1_cmd_ready             ),
  .i8_icb_cmd_sel                 (xbar_mg5_ro_to_sg1_cmd_sel               ),
  .i8_icb_cmd_read                (xbar_mg5_ro_to_sg1_cmd_read              ),
  .i8_icb_cmd_addr                (xbar_mg5_ro_to_sg1_cmd_addr   [  31:   0]),
  .i8_icb_cmd_wdata               (xbar_mg5_ro_to_sg1_cmd_wdata  [  63:   0]),
  .i8_icb_cmd_wmask               (xbar_mg5_ro_to_sg1_cmd_wmask  [   7:   0]),
  .i8_icb_cmd_size                (xbar_mg5_ro_to_sg1_cmd_size   [   2:   0]),
  .i8_icb_cmd_lock                (xbar_mg5_ro_to_sg1_cmd_lock              ),
  .i8_icb_cmd_excl                (xbar_mg5_ro_to_sg1_cmd_excl              ),
  .i8_icb_cmd_xlen                (xbar_mg5_ro_to_sg1_cmd_xlen   [   7:   0]),
  .i8_icb_cmd_xburst              (xbar_mg5_ro_to_sg1_cmd_xburst [   1:   0]),
  .i8_icb_cmd_modes               (xbar_mg5_ro_to_sg1_cmd_modes  [   1:   0]),
  .i8_icb_cmd_dmode               (xbar_mg5_ro_to_sg1_cmd_dmode             ),
  .i8_icb_cmd_attri               (xbar_mg5_ro_to_sg1_cmd_attri  [   2:   0]),
  .i8_icb_cmd_beat                (xbar_mg5_ro_to_sg1_cmd_beat   [   1:   0]),
  .i8_icb_cmd_usr                 (xbar_mg5_ro_to_sg1_cmd_usr    [   2:   0]),
  .i8_icb_rsp_ready               (xbar_mg5_ro_to_sg1_rsp_ready             ),
  .i8_icb_rsp_valid               (xbar_mg5_ro_to_sg1_rsp_valid             ),
  .i8_icb_rsp_err                 (xbar_mg5_ro_to_sg1_rsp_err               ),
  .i8_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg1_rsp_excl_ok            ),
  .i8_icb_rsp_rdata               (xbar_mg5_ro_to_sg1_rsp_rdata  [  63:   0]),
  .i8_icb_rsp_usr                 (xbar_mg5_ro_to_sg1_rsp_usr    [   2:   0]),
      .i9_icb_cmd_valid               (xbar_mg5_wo_to_sg1_cmd_valid             ),
  .i9_icb_cmd_ready               (xbar_mg5_wo_to_sg1_cmd_ready             ),
  .i9_icb_cmd_sel                 (xbar_mg5_wo_to_sg1_cmd_sel               ),
  .i9_icb_cmd_read                (xbar_mg5_wo_to_sg1_cmd_read              ),
  .i9_icb_cmd_addr                (xbar_mg5_wo_to_sg1_cmd_addr   [  31:   0]),
  .i9_icb_cmd_wdata               (xbar_mg5_wo_to_sg1_cmd_wdata  [  63:   0]),
  .i9_icb_cmd_wmask               (xbar_mg5_wo_to_sg1_cmd_wmask  [   7:   0]),
  .i9_icb_cmd_size                (xbar_mg5_wo_to_sg1_cmd_size   [   2:   0]),
  .i9_icb_cmd_lock                (xbar_mg5_wo_to_sg1_cmd_lock              ),
  .i9_icb_cmd_excl                (xbar_mg5_wo_to_sg1_cmd_excl              ),
  .i9_icb_cmd_xlen                (xbar_mg5_wo_to_sg1_cmd_xlen   [   7:   0]),
  .i9_icb_cmd_xburst              (xbar_mg5_wo_to_sg1_cmd_xburst [   1:   0]),
  .i9_icb_cmd_modes               (xbar_mg5_wo_to_sg1_cmd_modes  [   1:   0]),
  .i9_icb_cmd_dmode               (xbar_mg5_wo_to_sg1_cmd_dmode             ),
  .i9_icb_cmd_attri               (xbar_mg5_wo_to_sg1_cmd_attri  [   2:   0]),
  .i9_icb_cmd_beat                (xbar_mg5_wo_to_sg1_cmd_beat   [   1:   0]),
  .i9_icb_cmd_usr                 (xbar_mg5_wo_to_sg1_cmd_usr    [   2:   0]),
  .i9_icb_rsp_ready               (xbar_mg5_wo_to_sg1_rsp_ready             ),
  .i9_icb_rsp_valid               (xbar_mg5_wo_to_sg1_rsp_valid             ),
  .i9_icb_rsp_err                 (xbar_mg5_wo_to_sg1_rsp_err               ),
  .i9_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg1_rsp_excl_ok            ),
  .i9_icb_rsp_rdata               (xbar_mg5_wo_to_sg1_rsp_rdata  [  63:   0]),
  .i9_icb_rsp_usr                 (xbar_mg5_wo_to_sg1_rsp_usr    [   2:   0]),
      .i10_icb_cmd_valid              (xbar_mg6_ro_to_sg1_cmd_valid             ),
  .i10_icb_cmd_ready              (xbar_mg6_ro_to_sg1_cmd_ready             ),
  .i10_icb_cmd_sel                (xbar_mg6_ro_to_sg1_cmd_sel               ),
  .i10_icb_cmd_read               (xbar_mg6_ro_to_sg1_cmd_read              ),
  .i10_icb_cmd_addr               (xbar_mg6_ro_to_sg1_cmd_addr   [  31:   0]),
  .i10_icb_cmd_wdata              (xbar_mg6_ro_to_sg1_cmd_wdata  [  63:   0]),
  .i10_icb_cmd_wmask              (xbar_mg6_ro_to_sg1_cmd_wmask  [   7:   0]),
  .i10_icb_cmd_size               (xbar_mg6_ro_to_sg1_cmd_size   [   2:   0]),
  .i10_icb_cmd_lock               (xbar_mg6_ro_to_sg1_cmd_lock              ),
  .i10_icb_cmd_excl               (xbar_mg6_ro_to_sg1_cmd_excl              ),
  .i10_icb_cmd_xlen               (xbar_mg6_ro_to_sg1_cmd_xlen   [   7:   0]),
  .i10_icb_cmd_xburst             (xbar_mg6_ro_to_sg1_cmd_xburst [   1:   0]),
  .i10_icb_cmd_modes              (xbar_mg6_ro_to_sg1_cmd_modes  [   1:   0]),
  .i10_icb_cmd_dmode              (xbar_mg6_ro_to_sg1_cmd_dmode             ),
  .i10_icb_cmd_attri              (xbar_mg6_ro_to_sg1_cmd_attri  [   2:   0]),
  .i10_icb_cmd_beat               (xbar_mg6_ro_to_sg1_cmd_beat   [   1:   0]),
  .i10_icb_cmd_usr                (xbar_mg6_ro_to_sg1_cmd_usr    [   2:   0]),
  .i10_icb_rsp_ready              (xbar_mg6_ro_to_sg1_rsp_ready             ),
  .i10_icb_rsp_valid              (xbar_mg6_ro_to_sg1_rsp_valid             ),
  .i10_icb_rsp_err                (xbar_mg6_ro_to_sg1_rsp_err               ),
  .i10_icb_rsp_excl_ok            (xbar_mg6_ro_to_sg1_rsp_excl_ok            ),
  .i10_icb_rsp_rdata              (xbar_mg6_ro_to_sg1_rsp_rdata  [  63:   0]),
  .i10_icb_rsp_usr                (xbar_mg6_ro_to_sg1_rsp_usr    [   2:   0]),
      .i11_icb_cmd_valid              (xbar_mg6_wo_to_sg1_cmd_valid             ),
  .i11_icb_cmd_ready              (xbar_mg6_wo_to_sg1_cmd_ready             ),
  .i11_icb_cmd_sel                (xbar_mg6_wo_to_sg1_cmd_sel               ),
  .i11_icb_cmd_read               (xbar_mg6_wo_to_sg1_cmd_read              ),
  .i11_icb_cmd_addr               (xbar_mg6_wo_to_sg1_cmd_addr   [  31:   0]),
  .i11_icb_cmd_wdata              (xbar_mg6_wo_to_sg1_cmd_wdata  [  63:   0]),
  .i11_icb_cmd_wmask              (xbar_mg6_wo_to_sg1_cmd_wmask  [   7:   0]),
  .i11_icb_cmd_size               (xbar_mg6_wo_to_sg1_cmd_size   [   2:   0]),
  .i11_icb_cmd_lock               (xbar_mg6_wo_to_sg1_cmd_lock              ),
  .i11_icb_cmd_excl               (xbar_mg6_wo_to_sg1_cmd_excl              ),
  .i11_icb_cmd_xlen               (xbar_mg6_wo_to_sg1_cmd_xlen   [   7:   0]),
  .i11_icb_cmd_xburst             (xbar_mg6_wo_to_sg1_cmd_xburst [   1:   0]),
  .i11_icb_cmd_modes              (xbar_mg6_wo_to_sg1_cmd_modes  [   1:   0]),
  .i11_icb_cmd_dmode              (xbar_mg6_wo_to_sg1_cmd_dmode             ),
  .i11_icb_cmd_attri              (xbar_mg6_wo_to_sg1_cmd_attri  [   2:   0]),
  .i11_icb_cmd_beat               (xbar_mg6_wo_to_sg1_cmd_beat   [   1:   0]),
  .i11_icb_cmd_usr                (xbar_mg6_wo_to_sg1_cmd_usr    [   2:   0]),
  .i11_icb_rsp_ready              (xbar_mg6_wo_to_sg1_rsp_ready             ),
  .i11_icb_rsp_valid              (xbar_mg6_wo_to_sg1_rsp_valid             ),
  .i11_icb_rsp_err                (xbar_mg6_wo_to_sg1_rsp_err               ),
  .i11_icb_rsp_excl_ok            (xbar_mg6_wo_to_sg1_rsp_excl_ok            ),
  .i11_icb_rsp_rdata              (xbar_mg6_wo_to_sg1_rsp_rdata  [  63:   0]),
  .i11_icb_rsp_usr                (xbar_mg6_wo_to_sg1_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg2_rw_arbt_active;
   e603_subsys_xbar_slv2_rw_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (16  ),
      .ARBT_FIFO_OUTS_CNT_W(5),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg2_rw_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg2_rw_arbt_active),
      .o_icb_cmd_valid                (slv_grp_2_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (slv_grp_2_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (slv_grp_2_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (slv_grp_2_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (slv_grp_2_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_2_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_2_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_2_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_2_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (slv_grp_2_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (slv_grp_2_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_2_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_2_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_2_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (slv_grp_2_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_2_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_2_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_2_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (slv_grp_2_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (slv_grp_2_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (slv_grp_2_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (slv_grp_2_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_2_icb_rsp_usr         [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_ro_to_sg2_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_ro_to_sg2_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_ro_to_sg2_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_ro_to_sg2_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_ro_to_sg2_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_ro_to_sg2_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_ro_to_sg2_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_ro_to_sg2_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_ro_to_sg2_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_ro_to_sg2_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_ro_to_sg2_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_ro_to_sg2_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_ro_to_sg2_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_ro_to_sg2_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_ro_to_sg2_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_ro_to_sg2_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_ro_to_sg2_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_ro_to_sg2_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_ro_to_sg2_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_ro_to_sg2_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg2_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_ro_to_sg2_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_ro_to_sg2_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg0_wo_to_sg2_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg0_wo_to_sg2_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg0_wo_to_sg2_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg0_wo_to_sg2_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg0_wo_to_sg2_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg0_wo_to_sg2_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg0_wo_to_sg2_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg0_wo_to_sg2_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg0_wo_to_sg2_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg0_wo_to_sg2_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg0_wo_to_sg2_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg0_wo_to_sg2_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg0_wo_to_sg2_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg0_wo_to_sg2_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg0_wo_to_sg2_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg0_wo_to_sg2_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg0_wo_to_sg2_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg0_wo_to_sg2_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg0_wo_to_sg2_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg0_wo_to_sg2_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg2_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg0_wo_to_sg2_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg0_wo_to_sg2_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg1_ro_to_sg2_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg1_ro_to_sg2_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg1_ro_to_sg2_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg1_ro_to_sg2_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg1_ro_to_sg2_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg1_ro_to_sg2_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg1_ro_to_sg2_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg1_ro_to_sg2_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg1_ro_to_sg2_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg1_ro_to_sg2_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg1_ro_to_sg2_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg1_ro_to_sg2_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg1_ro_to_sg2_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg1_ro_to_sg2_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg1_ro_to_sg2_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg1_ro_to_sg2_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg1_ro_to_sg2_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg1_ro_to_sg2_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg1_ro_to_sg2_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg1_ro_to_sg2_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg2_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg1_ro_to_sg2_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg1_ro_to_sg2_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg2_wo_to_sg2_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg2_wo_to_sg2_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg2_wo_to_sg2_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg2_wo_to_sg2_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg2_wo_to_sg2_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg2_wo_to_sg2_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg2_wo_to_sg2_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg2_wo_to_sg2_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg2_wo_to_sg2_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg2_wo_to_sg2_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg2_wo_to_sg2_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg2_wo_to_sg2_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg2_wo_to_sg2_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg2_wo_to_sg2_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg2_wo_to_sg2_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg2_wo_to_sg2_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg2_wo_to_sg2_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg2_wo_to_sg2_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg2_wo_to_sg2_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg2_wo_to_sg2_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg2_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg2_wo_to_sg2_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg2_wo_to_sg2_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg3_ro_to_sg2_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg3_ro_to_sg2_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg3_ro_to_sg2_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg3_ro_to_sg2_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg3_ro_to_sg2_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg3_ro_to_sg2_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg3_ro_to_sg2_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg3_ro_to_sg2_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg3_ro_to_sg2_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg3_ro_to_sg2_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg3_ro_to_sg2_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg3_ro_to_sg2_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg3_ro_to_sg2_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg3_ro_to_sg2_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg3_ro_to_sg2_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg3_ro_to_sg2_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg3_ro_to_sg2_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg3_ro_to_sg2_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg3_ro_to_sg2_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg3_ro_to_sg2_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg2_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg3_ro_to_sg2_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg3_ro_to_sg2_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg3_wo_to_sg2_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg3_wo_to_sg2_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg3_wo_to_sg2_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg3_wo_to_sg2_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg3_wo_to_sg2_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg3_wo_to_sg2_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg3_wo_to_sg2_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg3_wo_to_sg2_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg3_wo_to_sg2_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg3_wo_to_sg2_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg3_wo_to_sg2_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg3_wo_to_sg2_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg3_wo_to_sg2_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg3_wo_to_sg2_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg3_wo_to_sg2_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg3_wo_to_sg2_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg3_wo_to_sg2_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg3_wo_to_sg2_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg3_wo_to_sg2_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg3_wo_to_sg2_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg2_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg3_wo_to_sg2_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg3_wo_to_sg2_rsp_usr    [   2:   0]),
      .i6_icb_cmd_valid               (xbar_mg4_ro_to_sg2_cmd_valid             ),
  .i6_icb_cmd_ready               (xbar_mg4_ro_to_sg2_cmd_ready             ),
  .i6_icb_cmd_sel                 (xbar_mg4_ro_to_sg2_cmd_sel               ),
  .i6_icb_cmd_read                (xbar_mg4_ro_to_sg2_cmd_read              ),
  .i6_icb_cmd_addr                (xbar_mg4_ro_to_sg2_cmd_addr   [  31:   0]),
  .i6_icb_cmd_wdata               (xbar_mg4_ro_to_sg2_cmd_wdata  [  63:   0]),
  .i6_icb_cmd_wmask               (xbar_mg4_ro_to_sg2_cmd_wmask  [   7:   0]),
  .i6_icb_cmd_size                (xbar_mg4_ro_to_sg2_cmd_size   [   2:   0]),
  .i6_icb_cmd_lock                (xbar_mg4_ro_to_sg2_cmd_lock              ),
  .i6_icb_cmd_excl                (xbar_mg4_ro_to_sg2_cmd_excl              ),
  .i6_icb_cmd_xlen                (xbar_mg4_ro_to_sg2_cmd_xlen   [   7:   0]),
  .i6_icb_cmd_xburst              (xbar_mg4_ro_to_sg2_cmd_xburst [   1:   0]),
  .i6_icb_cmd_modes               (xbar_mg4_ro_to_sg2_cmd_modes  [   1:   0]),
  .i6_icb_cmd_dmode               (xbar_mg4_ro_to_sg2_cmd_dmode             ),
  .i6_icb_cmd_attri               (xbar_mg4_ro_to_sg2_cmd_attri  [   2:   0]),
  .i6_icb_cmd_beat                (xbar_mg4_ro_to_sg2_cmd_beat   [   1:   0]),
  .i6_icb_cmd_usr                 (xbar_mg4_ro_to_sg2_cmd_usr    [   2:   0]),
  .i6_icb_rsp_ready               (xbar_mg4_ro_to_sg2_rsp_ready             ),
  .i6_icb_rsp_valid               (xbar_mg4_ro_to_sg2_rsp_valid             ),
  .i6_icb_rsp_err                 (xbar_mg4_ro_to_sg2_rsp_err               ),
  .i6_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg2_rsp_excl_ok            ),
  .i6_icb_rsp_rdata               (xbar_mg4_ro_to_sg2_rsp_rdata  [  63:   0]),
  .i6_icb_rsp_usr                 (xbar_mg4_ro_to_sg2_rsp_usr    [   2:   0]),
      .i7_icb_cmd_valid               (xbar_mg4_wo_to_sg2_cmd_valid             ),
  .i7_icb_cmd_ready               (xbar_mg4_wo_to_sg2_cmd_ready             ),
  .i7_icb_cmd_sel                 (xbar_mg4_wo_to_sg2_cmd_sel               ),
  .i7_icb_cmd_read                (xbar_mg4_wo_to_sg2_cmd_read              ),
  .i7_icb_cmd_addr                (xbar_mg4_wo_to_sg2_cmd_addr   [  31:   0]),
  .i7_icb_cmd_wdata               (xbar_mg4_wo_to_sg2_cmd_wdata  [  63:   0]),
  .i7_icb_cmd_wmask               (xbar_mg4_wo_to_sg2_cmd_wmask  [   7:   0]),
  .i7_icb_cmd_size                (xbar_mg4_wo_to_sg2_cmd_size   [   2:   0]),
  .i7_icb_cmd_lock                (xbar_mg4_wo_to_sg2_cmd_lock              ),
  .i7_icb_cmd_excl                (xbar_mg4_wo_to_sg2_cmd_excl              ),
  .i7_icb_cmd_xlen                (xbar_mg4_wo_to_sg2_cmd_xlen   [   7:   0]),
  .i7_icb_cmd_xburst              (xbar_mg4_wo_to_sg2_cmd_xburst [   1:   0]),
  .i7_icb_cmd_modes               (xbar_mg4_wo_to_sg2_cmd_modes  [   1:   0]),
  .i7_icb_cmd_dmode               (xbar_mg4_wo_to_sg2_cmd_dmode             ),
  .i7_icb_cmd_attri               (xbar_mg4_wo_to_sg2_cmd_attri  [   2:   0]),
  .i7_icb_cmd_beat                (xbar_mg4_wo_to_sg2_cmd_beat   [   1:   0]),
  .i7_icb_cmd_usr                 (xbar_mg4_wo_to_sg2_cmd_usr    [   2:   0]),
  .i7_icb_rsp_ready               (xbar_mg4_wo_to_sg2_rsp_ready             ),
  .i7_icb_rsp_valid               (xbar_mg4_wo_to_sg2_rsp_valid             ),
  .i7_icb_rsp_err                 (xbar_mg4_wo_to_sg2_rsp_err               ),
  .i7_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg2_rsp_excl_ok            ),
  .i7_icb_rsp_rdata               (xbar_mg4_wo_to_sg2_rsp_rdata  [  63:   0]),
  .i7_icb_rsp_usr                 (xbar_mg4_wo_to_sg2_rsp_usr    [   2:   0]),
      .i8_icb_cmd_valid               (xbar_mg5_ro_to_sg2_cmd_valid             ),
  .i8_icb_cmd_ready               (xbar_mg5_ro_to_sg2_cmd_ready             ),
  .i8_icb_cmd_sel                 (xbar_mg5_ro_to_sg2_cmd_sel               ),
  .i8_icb_cmd_read                (xbar_mg5_ro_to_sg2_cmd_read              ),
  .i8_icb_cmd_addr                (xbar_mg5_ro_to_sg2_cmd_addr   [  31:   0]),
  .i8_icb_cmd_wdata               (xbar_mg5_ro_to_sg2_cmd_wdata  [  63:   0]),
  .i8_icb_cmd_wmask               (xbar_mg5_ro_to_sg2_cmd_wmask  [   7:   0]),
  .i8_icb_cmd_size                (xbar_mg5_ro_to_sg2_cmd_size   [   2:   0]),
  .i8_icb_cmd_lock                (xbar_mg5_ro_to_sg2_cmd_lock              ),
  .i8_icb_cmd_excl                (xbar_mg5_ro_to_sg2_cmd_excl              ),
  .i8_icb_cmd_xlen                (xbar_mg5_ro_to_sg2_cmd_xlen   [   7:   0]),
  .i8_icb_cmd_xburst              (xbar_mg5_ro_to_sg2_cmd_xburst [   1:   0]),
  .i8_icb_cmd_modes               (xbar_mg5_ro_to_sg2_cmd_modes  [   1:   0]),
  .i8_icb_cmd_dmode               (xbar_mg5_ro_to_sg2_cmd_dmode             ),
  .i8_icb_cmd_attri               (xbar_mg5_ro_to_sg2_cmd_attri  [   2:   0]),
  .i8_icb_cmd_beat                (xbar_mg5_ro_to_sg2_cmd_beat   [   1:   0]),
  .i8_icb_cmd_usr                 (xbar_mg5_ro_to_sg2_cmd_usr    [   2:   0]),
  .i8_icb_rsp_ready               (xbar_mg5_ro_to_sg2_rsp_ready             ),
  .i8_icb_rsp_valid               (xbar_mg5_ro_to_sg2_rsp_valid             ),
  .i8_icb_rsp_err                 (xbar_mg5_ro_to_sg2_rsp_err               ),
  .i8_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg2_rsp_excl_ok            ),
  .i8_icb_rsp_rdata               (xbar_mg5_ro_to_sg2_rsp_rdata  [  63:   0]),
  .i8_icb_rsp_usr                 (xbar_mg5_ro_to_sg2_rsp_usr    [   2:   0]),
      .i9_icb_cmd_valid               (xbar_mg5_wo_to_sg2_cmd_valid             ),
  .i9_icb_cmd_ready               (xbar_mg5_wo_to_sg2_cmd_ready             ),
  .i9_icb_cmd_sel                 (xbar_mg5_wo_to_sg2_cmd_sel               ),
  .i9_icb_cmd_read                (xbar_mg5_wo_to_sg2_cmd_read              ),
  .i9_icb_cmd_addr                (xbar_mg5_wo_to_sg2_cmd_addr   [  31:   0]),
  .i9_icb_cmd_wdata               (xbar_mg5_wo_to_sg2_cmd_wdata  [  63:   0]),
  .i9_icb_cmd_wmask               (xbar_mg5_wo_to_sg2_cmd_wmask  [   7:   0]),
  .i9_icb_cmd_size                (xbar_mg5_wo_to_sg2_cmd_size   [   2:   0]),
  .i9_icb_cmd_lock                (xbar_mg5_wo_to_sg2_cmd_lock              ),
  .i9_icb_cmd_excl                (xbar_mg5_wo_to_sg2_cmd_excl              ),
  .i9_icb_cmd_xlen                (xbar_mg5_wo_to_sg2_cmd_xlen   [   7:   0]),
  .i9_icb_cmd_xburst              (xbar_mg5_wo_to_sg2_cmd_xburst [   1:   0]),
  .i9_icb_cmd_modes               (xbar_mg5_wo_to_sg2_cmd_modes  [   1:   0]),
  .i9_icb_cmd_dmode               (xbar_mg5_wo_to_sg2_cmd_dmode             ),
  .i9_icb_cmd_attri               (xbar_mg5_wo_to_sg2_cmd_attri  [   2:   0]),
  .i9_icb_cmd_beat                (xbar_mg5_wo_to_sg2_cmd_beat   [   1:   0]),
  .i9_icb_cmd_usr                 (xbar_mg5_wo_to_sg2_cmd_usr    [   2:   0]),
  .i9_icb_rsp_ready               (xbar_mg5_wo_to_sg2_rsp_ready             ),
  .i9_icb_rsp_valid               (xbar_mg5_wo_to_sg2_rsp_valid             ),
  .i9_icb_rsp_err                 (xbar_mg5_wo_to_sg2_rsp_err               ),
  .i9_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg2_rsp_excl_ok            ),
  .i9_icb_rsp_rdata               (xbar_mg5_wo_to_sg2_rsp_rdata  [  63:   0]),
  .i9_icb_rsp_usr                 (xbar_mg5_wo_to_sg2_rsp_usr    [   2:   0]),
      .i10_icb_cmd_valid              (xbar_mg6_ro_to_sg2_cmd_valid             ),
  .i10_icb_cmd_ready              (xbar_mg6_ro_to_sg2_cmd_ready             ),
  .i10_icb_cmd_sel                (xbar_mg6_ro_to_sg2_cmd_sel               ),
  .i10_icb_cmd_read               (xbar_mg6_ro_to_sg2_cmd_read              ),
  .i10_icb_cmd_addr               (xbar_mg6_ro_to_sg2_cmd_addr   [  31:   0]),
  .i10_icb_cmd_wdata              (xbar_mg6_ro_to_sg2_cmd_wdata  [  63:   0]),
  .i10_icb_cmd_wmask              (xbar_mg6_ro_to_sg2_cmd_wmask  [   7:   0]),
  .i10_icb_cmd_size               (xbar_mg6_ro_to_sg2_cmd_size   [   2:   0]),
  .i10_icb_cmd_lock               (xbar_mg6_ro_to_sg2_cmd_lock              ),
  .i10_icb_cmd_excl               (xbar_mg6_ro_to_sg2_cmd_excl              ),
  .i10_icb_cmd_xlen               (xbar_mg6_ro_to_sg2_cmd_xlen   [   7:   0]),
  .i10_icb_cmd_xburst             (xbar_mg6_ro_to_sg2_cmd_xburst [   1:   0]),
  .i10_icb_cmd_modes              (xbar_mg6_ro_to_sg2_cmd_modes  [   1:   0]),
  .i10_icb_cmd_dmode              (xbar_mg6_ro_to_sg2_cmd_dmode             ),
  .i10_icb_cmd_attri              (xbar_mg6_ro_to_sg2_cmd_attri  [   2:   0]),
  .i10_icb_cmd_beat               (xbar_mg6_ro_to_sg2_cmd_beat   [   1:   0]),
  .i10_icb_cmd_usr                (xbar_mg6_ro_to_sg2_cmd_usr    [   2:   0]),
  .i10_icb_rsp_ready              (xbar_mg6_ro_to_sg2_rsp_ready             ),
  .i10_icb_rsp_valid              (xbar_mg6_ro_to_sg2_rsp_valid             ),
  .i10_icb_rsp_err                (xbar_mg6_ro_to_sg2_rsp_err               ),
  .i10_icb_rsp_excl_ok            (xbar_mg6_ro_to_sg2_rsp_excl_ok            ),
  .i10_icb_rsp_rdata              (xbar_mg6_ro_to_sg2_rsp_rdata  [  63:   0]),
  .i10_icb_rsp_usr                (xbar_mg6_ro_to_sg2_rsp_usr    [   2:   0]),
      .i11_icb_cmd_valid              (xbar_mg6_wo_to_sg2_cmd_valid             ),
  .i11_icb_cmd_ready              (xbar_mg6_wo_to_sg2_cmd_ready             ),
  .i11_icb_cmd_sel                (xbar_mg6_wo_to_sg2_cmd_sel               ),
  .i11_icb_cmd_read               (xbar_mg6_wo_to_sg2_cmd_read              ),
  .i11_icb_cmd_addr               (xbar_mg6_wo_to_sg2_cmd_addr   [  31:   0]),
  .i11_icb_cmd_wdata              (xbar_mg6_wo_to_sg2_cmd_wdata  [  63:   0]),
  .i11_icb_cmd_wmask              (xbar_mg6_wo_to_sg2_cmd_wmask  [   7:   0]),
  .i11_icb_cmd_size               (xbar_mg6_wo_to_sg2_cmd_size   [   2:   0]),
  .i11_icb_cmd_lock               (xbar_mg6_wo_to_sg2_cmd_lock              ),
  .i11_icb_cmd_excl               (xbar_mg6_wo_to_sg2_cmd_excl              ),
  .i11_icb_cmd_xlen               (xbar_mg6_wo_to_sg2_cmd_xlen   [   7:   0]),
  .i11_icb_cmd_xburst             (xbar_mg6_wo_to_sg2_cmd_xburst [   1:   0]),
  .i11_icb_cmd_modes              (xbar_mg6_wo_to_sg2_cmd_modes  [   1:   0]),
  .i11_icb_cmd_dmode              (xbar_mg6_wo_to_sg2_cmd_dmode             ),
  .i11_icb_cmd_attri              (xbar_mg6_wo_to_sg2_cmd_attri  [   2:   0]),
  .i11_icb_cmd_beat               (xbar_mg6_wo_to_sg2_cmd_beat   [   1:   0]),
  .i11_icb_cmd_usr                (xbar_mg6_wo_to_sg2_cmd_usr    [   2:   0]),
  .i11_icb_rsp_ready              (xbar_mg6_wo_to_sg2_rsp_ready             ),
  .i11_icb_rsp_valid              (xbar_mg6_wo_to_sg2_rsp_valid             ),
  .i11_icb_rsp_err                (xbar_mg6_wo_to_sg2_rsp_err               ),
  .i11_icb_rsp_excl_ok            (xbar_mg6_wo_to_sg2_rsp_excl_ok            ),
  .i11_icb_rsp_rdata              (xbar_mg6_wo_to_sg2_rsp_rdata  [  63:   0]),
  .i11_icb_rsp_usr                (xbar_mg6_wo_to_sg2_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg3_rw_arbt_active;
   e603_subsys_xbar_slv3_rw_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (16  ),
      .ARBT_FIFO_OUTS_CNT_W(5),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg3_rw_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg3_rw_arbt_active),
      .o_icb_cmd_valid                (slv_grp_3_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (slv_grp_3_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (slv_grp_3_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (slv_grp_3_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (slv_grp_3_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_3_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_3_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_3_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_3_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (slv_grp_3_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (slv_grp_3_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_3_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_3_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_3_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (slv_grp_3_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_3_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_3_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_3_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (slv_grp_3_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (slv_grp_3_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (slv_grp_3_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (slv_grp_3_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_3_icb_rsp_usr         [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_ro_to_sg3_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_ro_to_sg3_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_ro_to_sg3_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_ro_to_sg3_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_ro_to_sg3_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_ro_to_sg3_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_ro_to_sg3_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_ro_to_sg3_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_ro_to_sg3_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_ro_to_sg3_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_ro_to_sg3_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_ro_to_sg3_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_ro_to_sg3_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_ro_to_sg3_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_ro_to_sg3_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_ro_to_sg3_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_ro_to_sg3_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_ro_to_sg3_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_ro_to_sg3_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_ro_to_sg3_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg3_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_ro_to_sg3_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_ro_to_sg3_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg0_wo_to_sg3_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg0_wo_to_sg3_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg0_wo_to_sg3_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg0_wo_to_sg3_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg0_wo_to_sg3_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg0_wo_to_sg3_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg0_wo_to_sg3_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg0_wo_to_sg3_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg0_wo_to_sg3_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg0_wo_to_sg3_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg0_wo_to_sg3_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg0_wo_to_sg3_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg0_wo_to_sg3_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg0_wo_to_sg3_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg0_wo_to_sg3_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg0_wo_to_sg3_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg0_wo_to_sg3_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg0_wo_to_sg3_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg0_wo_to_sg3_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg0_wo_to_sg3_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg3_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg0_wo_to_sg3_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg0_wo_to_sg3_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg1_ro_to_sg3_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg1_ro_to_sg3_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg1_ro_to_sg3_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg1_ro_to_sg3_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg1_ro_to_sg3_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg1_ro_to_sg3_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg1_ro_to_sg3_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg1_ro_to_sg3_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg1_ro_to_sg3_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg1_ro_to_sg3_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg1_ro_to_sg3_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg1_ro_to_sg3_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg1_ro_to_sg3_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg1_ro_to_sg3_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg1_ro_to_sg3_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg1_ro_to_sg3_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg1_ro_to_sg3_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg1_ro_to_sg3_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg1_ro_to_sg3_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg1_ro_to_sg3_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg3_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg1_ro_to_sg3_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg1_ro_to_sg3_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg2_wo_to_sg3_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg2_wo_to_sg3_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg2_wo_to_sg3_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg2_wo_to_sg3_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg2_wo_to_sg3_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg2_wo_to_sg3_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg2_wo_to_sg3_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg2_wo_to_sg3_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg2_wo_to_sg3_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg2_wo_to_sg3_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg2_wo_to_sg3_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg2_wo_to_sg3_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg2_wo_to_sg3_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg2_wo_to_sg3_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg2_wo_to_sg3_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg2_wo_to_sg3_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg2_wo_to_sg3_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg2_wo_to_sg3_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg2_wo_to_sg3_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg2_wo_to_sg3_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg3_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg2_wo_to_sg3_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg2_wo_to_sg3_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg3_ro_to_sg3_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg3_ro_to_sg3_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg3_ro_to_sg3_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg3_ro_to_sg3_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg3_ro_to_sg3_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg3_ro_to_sg3_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg3_ro_to_sg3_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg3_ro_to_sg3_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg3_ro_to_sg3_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg3_ro_to_sg3_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg3_ro_to_sg3_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg3_ro_to_sg3_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg3_ro_to_sg3_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg3_ro_to_sg3_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg3_ro_to_sg3_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg3_ro_to_sg3_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg3_ro_to_sg3_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg3_ro_to_sg3_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg3_ro_to_sg3_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg3_ro_to_sg3_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg3_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg3_ro_to_sg3_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg3_ro_to_sg3_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg3_wo_to_sg3_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg3_wo_to_sg3_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg3_wo_to_sg3_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg3_wo_to_sg3_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg3_wo_to_sg3_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg3_wo_to_sg3_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg3_wo_to_sg3_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg3_wo_to_sg3_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg3_wo_to_sg3_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg3_wo_to_sg3_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg3_wo_to_sg3_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg3_wo_to_sg3_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg3_wo_to_sg3_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg3_wo_to_sg3_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg3_wo_to_sg3_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg3_wo_to_sg3_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg3_wo_to_sg3_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg3_wo_to_sg3_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg3_wo_to_sg3_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg3_wo_to_sg3_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg3_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg3_wo_to_sg3_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg3_wo_to_sg3_rsp_usr    [   2:   0]),
      .i6_icb_cmd_valid               (xbar_mg4_ro_to_sg3_cmd_valid             ),
  .i6_icb_cmd_ready               (xbar_mg4_ro_to_sg3_cmd_ready             ),
  .i6_icb_cmd_sel                 (xbar_mg4_ro_to_sg3_cmd_sel               ),
  .i6_icb_cmd_read                (xbar_mg4_ro_to_sg3_cmd_read              ),
  .i6_icb_cmd_addr                (xbar_mg4_ro_to_sg3_cmd_addr   [  31:   0]),
  .i6_icb_cmd_wdata               (xbar_mg4_ro_to_sg3_cmd_wdata  [  63:   0]),
  .i6_icb_cmd_wmask               (xbar_mg4_ro_to_sg3_cmd_wmask  [   7:   0]),
  .i6_icb_cmd_size                (xbar_mg4_ro_to_sg3_cmd_size   [   2:   0]),
  .i6_icb_cmd_lock                (xbar_mg4_ro_to_sg3_cmd_lock              ),
  .i6_icb_cmd_excl                (xbar_mg4_ro_to_sg3_cmd_excl              ),
  .i6_icb_cmd_xlen                (xbar_mg4_ro_to_sg3_cmd_xlen   [   7:   0]),
  .i6_icb_cmd_xburst              (xbar_mg4_ro_to_sg3_cmd_xburst [   1:   0]),
  .i6_icb_cmd_modes               (xbar_mg4_ro_to_sg3_cmd_modes  [   1:   0]),
  .i6_icb_cmd_dmode               (xbar_mg4_ro_to_sg3_cmd_dmode             ),
  .i6_icb_cmd_attri               (xbar_mg4_ro_to_sg3_cmd_attri  [   2:   0]),
  .i6_icb_cmd_beat                (xbar_mg4_ro_to_sg3_cmd_beat   [   1:   0]),
  .i6_icb_cmd_usr                 (xbar_mg4_ro_to_sg3_cmd_usr    [   2:   0]),
  .i6_icb_rsp_ready               (xbar_mg4_ro_to_sg3_rsp_ready             ),
  .i6_icb_rsp_valid               (xbar_mg4_ro_to_sg3_rsp_valid             ),
  .i6_icb_rsp_err                 (xbar_mg4_ro_to_sg3_rsp_err               ),
  .i6_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg3_rsp_excl_ok            ),
  .i6_icb_rsp_rdata               (xbar_mg4_ro_to_sg3_rsp_rdata  [  63:   0]),
  .i6_icb_rsp_usr                 (xbar_mg4_ro_to_sg3_rsp_usr    [   2:   0]),
      .i7_icb_cmd_valid               (xbar_mg4_wo_to_sg3_cmd_valid             ),
  .i7_icb_cmd_ready               (xbar_mg4_wo_to_sg3_cmd_ready             ),
  .i7_icb_cmd_sel                 (xbar_mg4_wo_to_sg3_cmd_sel               ),
  .i7_icb_cmd_read                (xbar_mg4_wo_to_sg3_cmd_read              ),
  .i7_icb_cmd_addr                (xbar_mg4_wo_to_sg3_cmd_addr   [  31:   0]),
  .i7_icb_cmd_wdata               (xbar_mg4_wo_to_sg3_cmd_wdata  [  63:   0]),
  .i7_icb_cmd_wmask               (xbar_mg4_wo_to_sg3_cmd_wmask  [   7:   0]),
  .i7_icb_cmd_size                (xbar_mg4_wo_to_sg3_cmd_size   [   2:   0]),
  .i7_icb_cmd_lock                (xbar_mg4_wo_to_sg3_cmd_lock              ),
  .i7_icb_cmd_excl                (xbar_mg4_wo_to_sg3_cmd_excl              ),
  .i7_icb_cmd_xlen                (xbar_mg4_wo_to_sg3_cmd_xlen   [   7:   0]),
  .i7_icb_cmd_xburst              (xbar_mg4_wo_to_sg3_cmd_xburst [   1:   0]),
  .i7_icb_cmd_modes               (xbar_mg4_wo_to_sg3_cmd_modes  [   1:   0]),
  .i7_icb_cmd_dmode               (xbar_mg4_wo_to_sg3_cmd_dmode             ),
  .i7_icb_cmd_attri               (xbar_mg4_wo_to_sg3_cmd_attri  [   2:   0]),
  .i7_icb_cmd_beat                (xbar_mg4_wo_to_sg3_cmd_beat   [   1:   0]),
  .i7_icb_cmd_usr                 (xbar_mg4_wo_to_sg3_cmd_usr    [   2:   0]),
  .i7_icb_rsp_ready               (xbar_mg4_wo_to_sg3_rsp_ready             ),
  .i7_icb_rsp_valid               (xbar_mg4_wo_to_sg3_rsp_valid             ),
  .i7_icb_rsp_err                 (xbar_mg4_wo_to_sg3_rsp_err               ),
  .i7_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg3_rsp_excl_ok            ),
  .i7_icb_rsp_rdata               (xbar_mg4_wo_to_sg3_rsp_rdata  [  63:   0]),
  .i7_icb_rsp_usr                 (xbar_mg4_wo_to_sg3_rsp_usr    [   2:   0]),
      .i8_icb_cmd_valid               (xbar_mg5_ro_to_sg3_cmd_valid             ),
  .i8_icb_cmd_ready               (xbar_mg5_ro_to_sg3_cmd_ready             ),
  .i8_icb_cmd_sel                 (xbar_mg5_ro_to_sg3_cmd_sel               ),
  .i8_icb_cmd_read                (xbar_mg5_ro_to_sg3_cmd_read              ),
  .i8_icb_cmd_addr                (xbar_mg5_ro_to_sg3_cmd_addr   [  31:   0]),
  .i8_icb_cmd_wdata               (xbar_mg5_ro_to_sg3_cmd_wdata  [  63:   0]),
  .i8_icb_cmd_wmask               (xbar_mg5_ro_to_sg3_cmd_wmask  [   7:   0]),
  .i8_icb_cmd_size                (xbar_mg5_ro_to_sg3_cmd_size   [   2:   0]),
  .i8_icb_cmd_lock                (xbar_mg5_ro_to_sg3_cmd_lock              ),
  .i8_icb_cmd_excl                (xbar_mg5_ro_to_sg3_cmd_excl              ),
  .i8_icb_cmd_xlen                (xbar_mg5_ro_to_sg3_cmd_xlen   [   7:   0]),
  .i8_icb_cmd_xburst              (xbar_mg5_ro_to_sg3_cmd_xburst [   1:   0]),
  .i8_icb_cmd_modes               (xbar_mg5_ro_to_sg3_cmd_modes  [   1:   0]),
  .i8_icb_cmd_dmode               (xbar_mg5_ro_to_sg3_cmd_dmode             ),
  .i8_icb_cmd_attri               (xbar_mg5_ro_to_sg3_cmd_attri  [   2:   0]),
  .i8_icb_cmd_beat                (xbar_mg5_ro_to_sg3_cmd_beat   [   1:   0]),
  .i8_icb_cmd_usr                 (xbar_mg5_ro_to_sg3_cmd_usr    [   2:   0]),
  .i8_icb_rsp_ready               (xbar_mg5_ro_to_sg3_rsp_ready             ),
  .i8_icb_rsp_valid               (xbar_mg5_ro_to_sg3_rsp_valid             ),
  .i8_icb_rsp_err                 (xbar_mg5_ro_to_sg3_rsp_err               ),
  .i8_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg3_rsp_excl_ok            ),
  .i8_icb_rsp_rdata               (xbar_mg5_ro_to_sg3_rsp_rdata  [  63:   0]),
  .i8_icb_rsp_usr                 (xbar_mg5_ro_to_sg3_rsp_usr    [   2:   0]),
      .i9_icb_cmd_valid               (xbar_mg5_wo_to_sg3_cmd_valid             ),
  .i9_icb_cmd_ready               (xbar_mg5_wo_to_sg3_cmd_ready             ),
  .i9_icb_cmd_sel                 (xbar_mg5_wo_to_sg3_cmd_sel               ),
  .i9_icb_cmd_read                (xbar_mg5_wo_to_sg3_cmd_read              ),
  .i9_icb_cmd_addr                (xbar_mg5_wo_to_sg3_cmd_addr   [  31:   0]),
  .i9_icb_cmd_wdata               (xbar_mg5_wo_to_sg3_cmd_wdata  [  63:   0]),
  .i9_icb_cmd_wmask               (xbar_mg5_wo_to_sg3_cmd_wmask  [   7:   0]),
  .i9_icb_cmd_size                (xbar_mg5_wo_to_sg3_cmd_size   [   2:   0]),
  .i9_icb_cmd_lock                (xbar_mg5_wo_to_sg3_cmd_lock              ),
  .i9_icb_cmd_excl                (xbar_mg5_wo_to_sg3_cmd_excl              ),
  .i9_icb_cmd_xlen                (xbar_mg5_wo_to_sg3_cmd_xlen   [   7:   0]),
  .i9_icb_cmd_xburst              (xbar_mg5_wo_to_sg3_cmd_xburst [   1:   0]),
  .i9_icb_cmd_modes               (xbar_mg5_wo_to_sg3_cmd_modes  [   1:   0]),
  .i9_icb_cmd_dmode               (xbar_mg5_wo_to_sg3_cmd_dmode             ),
  .i9_icb_cmd_attri               (xbar_mg5_wo_to_sg3_cmd_attri  [   2:   0]),
  .i9_icb_cmd_beat                (xbar_mg5_wo_to_sg3_cmd_beat   [   1:   0]),
  .i9_icb_cmd_usr                 (xbar_mg5_wo_to_sg3_cmd_usr    [   2:   0]),
  .i9_icb_rsp_ready               (xbar_mg5_wo_to_sg3_rsp_ready             ),
  .i9_icb_rsp_valid               (xbar_mg5_wo_to_sg3_rsp_valid             ),
  .i9_icb_rsp_err                 (xbar_mg5_wo_to_sg3_rsp_err               ),
  .i9_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg3_rsp_excl_ok            ),
  .i9_icb_rsp_rdata               (xbar_mg5_wo_to_sg3_rsp_rdata  [  63:   0]),
  .i9_icb_rsp_usr                 (xbar_mg5_wo_to_sg3_rsp_usr    [   2:   0]),
      .i10_icb_cmd_valid              (xbar_mg6_ro_to_sg3_cmd_valid             ),
  .i10_icb_cmd_ready              (xbar_mg6_ro_to_sg3_cmd_ready             ),
  .i10_icb_cmd_sel                (xbar_mg6_ro_to_sg3_cmd_sel               ),
  .i10_icb_cmd_read               (xbar_mg6_ro_to_sg3_cmd_read              ),
  .i10_icb_cmd_addr               (xbar_mg6_ro_to_sg3_cmd_addr   [  31:   0]),
  .i10_icb_cmd_wdata              (xbar_mg6_ro_to_sg3_cmd_wdata  [  63:   0]),
  .i10_icb_cmd_wmask              (xbar_mg6_ro_to_sg3_cmd_wmask  [   7:   0]),
  .i10_icb_cmd_size               (xbar_mg6_ro_to_sg3_cmd_size   [   2:   0]),
  .i10_icb_cmd_lock               (xbar_mg6_ro_to_sg3_cmd_lock              ),
  .i10_icb_cmd_excl               (xbar_mg6_ro_to_sg3_cmd_excl              ),
  .i10_icb_cmd_xlen               (xbar_mg6_ro_to_sg3_cmd_xlen   [   7:   0]),
  .i10_icb_cmd_xburst             (xbar_mg6_ro_to_sg3_cmd_xburst [   1:   0]),
  .i10_icb_cmd_modes              (xbar_mg6_ro_to_sg3_cmd_modes  [   1:   0]),
  .i10_icb_cmd_dmode              (xbar_mg6_ro_to_sg3_cmd_dmode             ),
  .i10_icb_cmd_attri              (xbar_mg6_ro_to_sg3_cmd_attri  [   2:   0]),
  .i10_icb_cmd_beat               (xbar_mg6_ro_to_sg3_cmd_beat   [   1:   0]),
  .i10_icb_cmd_usr                (xbar_mg6_ro_to_sg3_cmd_usr    [   2:   0]),
  .i10_icb_rsp_ready              (xbar_mg6_ro_to_sg3_rsp_ready             ),
  .i10_icb_rsp_valid              (xbar_mg6_ro_to_sg3_rsp_valid             ),
  .i10_icb_rsp_err                (xbar_mg6_ro_to_sg3_rsp_err               ),
  .i10_icb_rsp_excl_ok            (xbar_mg6_ro_to_sg3_rsp_excl_ok            ),
  .i10_icb_rsp_rdata              (xbar_mg6_ro_to_sg3_rsp_rdata  [  63:   0]),
  .i10_icb_rsp_usr                (xbar_mg6_ro_to_sg3_rsp_usr    [   2:   0]),
      .i11_icb_cmd_valid              (xbar_mg6_wo_to_sg3_cmd_valid             ),
  .i11_icb_cmd_ready              (xbar_mg6_wo_to_sg3_cmd_ready             ),
  .i11_icb_cmd_sel                (xbar_mg6_wo_to_sg3_cmd_sel               ),
  .i11_icb_cmd_read               (xbar_mg6_wo_to_sg3_cmd_read              ),
  .i11_icb_cmd_addr               (xbar_mg6_wo_to_sg3_cmd_addr   [  31:   0]),
  .i11_icb_cmd_wdata              (xbar_mg6_wo_to_sg3_cmd_wdata  [  63:   0]),
  .i11_icb_cmd_wmask              (xbar_mg6_wo_to_sg3_cmd_wmask  [   7:   0]),
  .i11_icb_cmd_size               (xbar_mg6_wo_to_sg3_cmd_size   [   2:   0]),
  .i11_icb_cmd_lock               (xbar_mg6_wo_to_sg3_cmd_lock              ),
  .i11_icb_cmd_excl               (xbar_mg6_wo_to_sg3_cmd_excl              ),
  .i11_icb_cmd_xlen               (xbar_mg6_wo_to_sg3_cmd_xlen   [   7:   0]),
  .i11_icb_cmd_xburst             (xbar_mg6_wo_to_sg3_cmd_xburst [   1:   0]),
  .i11_icb_cmd_modes              (xbar_mg6_wo_to_sg3_cmd_modes  [   1:   0]),
  .i11_icb_cmd_dmode              (xbar_mg6_wo_to_sg3_cmd_dmode             ),
  .i11_icb_cmd_attri              (xbar_mg6_wo_to_sg3_cmd_attri  [   2:   0]),
  .i11_icb_cmd_beat               (xbar_mg6_wo_to_sg3_cmd_beat   [   1:   0]),
  .i11_icb_cmd_usr                (xbar_mg6_wo_to_sg3_cmd_usr    [   2:   0]),
  .i11_icb_rsp_ready              (xbar_mg6_wo_to_sg3_rsp_ready             ),
  .i11_icb_rsp_valid              (xbar_mg6_wo_to_sg3_rsp_valid             ),
  .i11_icb_rsp_err                (xbar_mg6_wo_to_sg3_rsp_err               ),
  .i11_icb_rsp_excl_ok            (xbar_mg6_wo_to_sg3_rsp_excl_ok            ),
  .i11_icb_rsp_rdata              (xbar_mg6_wo_to_sg3_rsp_rdata  [  63:   0]),
  .i11_icb_rsp_usr                (xbar_mg6_wo_to_sg3_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg4_rw_arbt_active;
   e603_subsys_xbar_slv4_rw_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (16  ),
      .ARBT_FIFO_OUTS_CNT_W(5),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg4_rw_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg4_rw_arbt_active),
      .o_icb_cmd_valid                (slv_grp_4_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (slv_grp_4_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (slv_grp_4_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (slv_grp_4_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (slv_grp_4_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_4_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_4_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_4_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_4_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (slv_grp_4_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (slv_grp_4_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_4_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_4_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_4_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (slv_grp_4_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_4_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_4_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_4_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (slv_grp_4_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (slv_grp_4_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (slv_grp_4_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (slv_grp_4_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_4_icb_rsp_usr         [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_ro_to_sg4_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_ro_to_sg4_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_ro_to_sg4_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_ro_to_sg4_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_ro_to_sg4_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_ro_to_sg4_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_ro_to_sg4_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_ro_to_sg4_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_ro_to_sg4_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_ro_to_sg4_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_ro_to_sg4_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_ro_to_sg4_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_ro_to_sg4_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_ro_to_sg4_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_ro_to_sg4_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_ro_to_sg4_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_ro_to_sg4_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_ro_to_sg4_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_ro_to_sg4_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_ro_to_sg4_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg4_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_ro_to_sg4_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_ro_to_sg4_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg0_wo_to_sg4_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg0_wo_to_sg4_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg0_wo_to_sg4_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg0_wo_to_sg4_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg0_wo_to_sg4_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg0_wo_to_sg4_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg0_wo_to_sg4_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg0_wo_to_sg4_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg0_wo_to_sg4_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg0_wo_to_sg4_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg0_wo_to_sg4_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg0_wo_to_sg4_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg0_wo_to_sg4_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg0_wo_to_sg4_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg0_wo_to_sg4_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg0_wo_to_sg4_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg0_wo_to_sg4_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg0_wo_to_sg4_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg0_wo_to_sg4_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg0_wo_to_sg4_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg4_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg0_wo_to_sg4_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg0_wo_to_sg4_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg1_ro_to_sg4_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg1_ro_to_sg4_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg1_ro_to_sg4_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg1_ro_to_sg4_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg1_ro_to_sg4_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg1_ro_to_sg4_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg1_ro_to_sg4_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg1_ro_to_sg4_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg1_ro_to_sg4_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg1_ro_to_sg4_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg1_ro_to_sg4_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg1_ro_to_sg4_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg1_ro_to_sg4_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg1_ro_to_sg4_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg1_ro_to_sg4_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg1_ro_to_sg4_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg1_ro_to_sg4_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg1_ro_to_sg4_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg1_ro_to_sg4_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg1_ro_to_sg4_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg4_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg1_ro_to_sg4_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg1_ro_to_sg4_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg2_wo_to_sg4_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg2_wo_to_sg4_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg2_wo_to_sg4_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg2_wo_to_sg4_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg2_wo_to_sg4_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg2_wo_to_sg4_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg2_wo_to_sg4_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg2_wo_to_sg4_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg2_wo_to_sg4_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg2_wo_to_sg4_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg2_wo_to_sg4_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg2_wo_to_sg4_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg2_wo_to_sg4_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg2_wo_to_sg4_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg2_wo_to_sg4_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg2_wo_to_sg4_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg2_wo_to_sg4_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg2_wo_to_sg4_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg2_wo_to_sg4_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg2_wo_to_sg4_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg4_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg2_wo_to_sg4_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg2_wo_to_sg4_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg3_ro_to_sg4_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg3_ro_to_sg4_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg3_ro_to_sg4_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg3_ro_to_sg4_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg3_ro_to_sg4_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg3_ro_to_sg4_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg3_ro_to_sg4_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg3_ro_to_sg4_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg3_ro_to_sg4_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg3_ro_to_sg4_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg3_ro_to_sg4_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg3_ro_to_sg4_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg3_ro_to_sg4_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg3_ro_to_sg4_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg3_ro_to_sg4_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg3_ro_to_sg4_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg3_ro_to_sg4_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg3_ro_to_sg4_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg3_ro_to_sg4_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg3_ro_to_sg4_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg4_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg3_ro_to_sg4_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg3_ro_to_sg4_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg3_wo_to_sg4_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg3_wo_to_sg4_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg3_wo_to_sg4_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg3_wo_to_sg4_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg3_wo_to_sg4_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg3_wo_to_sg4_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg3_wo_to_sg4_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg3_wo_to_sg4_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg3_wo_to_sg4_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg3_wo_to_sg4_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg3_wo_to_sg4_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg3_wo_to_sg4_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg3_wo_to_sg4_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg3_wo_to_sg4_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg3_wo_to_sg4_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg3_wo_to_sg4_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg3_wo_to_sg4_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg3_wo_to_sg4_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg3_wo_to_sg4_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg3_wo_to_sg4_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg4_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg3_wo_to_sg4_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg3_wo_to_sg4_rsp_usr    [   2:   0]),
      .i6_icb_cmd_valid               (xbar_mg4_ro_to_sg4_cmd_valid             ),
  .i6_icb_cmd_ready               (xbar_mg4_ro_to_sg4_cmd_ready             ),
  .i6_icb_cmd_sel                 (xbar_mg4_ro_to_sg4_cmd_sel               ),
  .i6_icb_cmd_read                (xbar_mg4_ro_to_sg4_cmd_read              ),
  .i6_icb_cmd_addr                (xbar_mg4_ro_to_sg4_cmd_addr   [  31:   0]),
  .i6_icb_cmd_wdata               (xbar_mg4_ro_to_sg4_cmd_wdata  [  63:   0]),
  .i6_icb_cmd_wmask               (xbar_mg4_ro_to_sg4_cmd_wmask  [   7:   0]),
  .i6_icb_cmd_size                (xbar_mg4_ro_to_sg4_cmd_size   [   2:   0]),
  .i6_icb_cmd_lock                (xbar_mg4_ro_to_sg4_cmd_lock              ),
  .i6_icb_cmd_excl                (xbar_mg4_ro_to_sg4_cmd_excl              ),
  .i6_icb_cmd_xlen                (xbar_mg4_ro_to_sg4_cmd_xlen   [   7:   0]),
  .i6_icb_cmd_xburst              (xbar_mg4_ro_to_sg4_cmd_xburst [   1:   0]),
  .i6_icb_cmd_modes               (xbar_mg4_ro_to_sg4_cmd_modes  [   1:   0]),
  .i6_icb_cmd_dmode               (xbar_mg4_ro_to_sg4_cmd_dmode             ),
  .i6_icb_cmd_attri               (xbar_mg4_ro_to_sg4_cmd_attri  [   2:   0]),
  .i6_icb_cmd_beat                (xbar_mg4_ro_to_sg4_cmd_beat   [   1:   0]),
  .i6_icb_cmd_usr                 (xbar_mg4_ro_to_sg4_cmd_usr    [   2:   0]),
  .i6_icb_rsp_ready               (xbar_mg4_ro_to_sg4_rsp_ready             ),
  .i6_icb_rsp_valid               (xbar_mg4_ro_to_sg4_rsp_valid             ),
  .i6_icb_rsp_err                 (xbar_mg4_ro_to_sg4_rsp_err               ),
  .i6_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg4_rsp_excl_ok            ),
  .i6_icb_rsp_rdata               (xbar_mg4_ro_to_sg4_rsp_rdata  [  63:   0]),
  .i6_icb_rsp_usr                 (xbar_mg4_ro_to_sg4_rsp_usr    [   2:   0]),
      .i7_icb_cmd_valid               (xbar_mg4_wo_to_sg4_cmd_valid             ),
  .i7_icb_cmd_ready               (xbar_mg4_wo_to_sg4_cmd_ready             ),
  .i7_icb_cmd_sel                 (xbar_mg4_wo_to_sg4_cmd_sel               ),
  .i7_icb_cmd_read                (xbar_mg4_wo_to_sg4_cmd_read              ),
  .i7_icb_cmd_addr                (xbar_mg4_wo_to_sg4_cmd_addr   [  31:   0]),
  .i7_icb_cmd_wdata               (xbar_mg4_wo_to_sg4_cmd_wdata  [  63:   0]),
  .i7_icb_cmd_wmask               (xbar_mg4_wo_to_sg4_cmd_wmask  [   7:   0]),
  .i7_icb_cmd_size                (xbar_mg4_wo_to_sg4_cmd_size   [   2:   0]),
  .i7_icb_cmd_lock                (xbar_mg4_wo_to_sg4_cmd_lock              ),
  .i7_icb_cmd_excl                (xbar_mg4_wo_to_sg4_cmd_excl              ),
  .i7_icb_cmd_xlen                (xbar_mg4_wo_to_sg4_cmd_xlen   [   7:   0]),
  .i7_icb_cmd_xburst              (xbar_mg4_wo_to_sg4_cmd_xburst [   1:   0]),
  .i7_icb_cmd_modes               (xbar_mg4_wo_to_sg4_cmd_modes  [   1:   0]),
  .i7_icb_cmd_dmode               (xbar_mg4_wo_to_sg4_cmd_dmode             ),
  .i7_icb_cmd_attri               (xbar_mg4_wo_to_sg4_cmd_attri  [   2:   0]),
  .i7_icb_cmd_beat                (xbar_mg4_wo_to_sg4_cmd_beat   [   1:   0]),
  .i7_icb_cmd_usr                 (xbar_mg4_wo_to_sg4_cmd_usr    [   2:   0]),
  .i7_icb_rsp_ready               (xbar_mg4_wo_to_sg4_rsp_ready             ),
  .i7_icb_rsp_valid               (xbar_mg4_wo_to_sg4_rsp_valid             ),
  .i7_icb_rsp_err                 (xbar_mg4_wo_to_sg4_rsp_err               ),
  .i7_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg4_rsp_excl_ok            ),
  .i7_icb_rsp_rdata               (xbar_mg4_wo_to_sg4_rsp_rdata  [  63:   0]),
  .i7_icb_rsp_usr                 (xbar_mg4_wo_to_sg4_rsp_usr    [   2:   0]),
      .i8_icb_cmd_valid               (xbar_mg5_ro_to_sg4_cmd_valid             ),
  .i8_icb_cmd_ready               (xbar_mg5_ro_to_sg4_cmd_ready             ),
  .i8_icb_cmd_sel                 (xbar_mg5_ro_to_sg4_cmd_sel               ),
  .i8_icb_cmd_read                (xbar_mg5_ro_to_sg4_cmd_read              ),
  .i8_icb_cmd_addr                (xbar_mg5_ro_to_sg4_cmd_addr   [  31:   0]),
  .i8_icb_cmd_wdata               (xbar_mg5_ro_to_sg4_cmd_wdata  [  63:   0]),
  .i8_icb_cmd_wmask               (xbar_mg5_ro_to_sg4_cmd_wmask  [   7:   0]),
  .i8_icb_cmd_size                (xbar_mg5_ro_to_sg4_cmd_size   [   2:   0]),
  .i8_icb_cmd_lock                (xbar_mg5_ro_to_sg4_cmd_lock              ),
  .i8_icb_cmd_excl                (xbar_mg5_ro_to_sg4_cmd_excl              ),
  .i8_icb_cmd_xlen                (xbar_mg5_ro_to_sg4_cmd_xlen   [   7:   0]),
  .i8_icb_cmd_xburst              (xbar_mg5_ro_to_sg4_cmd_xburst [   1:   0]),
  .i8_icb_cmd_modes               (xbar_mg5_ro_to_sg4_cmd_modes  [   1:   0]),
  .i8_icb_cmd_dmode               (xbar_mg5_ro_to_sg4_cmd_dmode             ),
  .i8_icb_cmd_attri               (xbar_mg5_ro_to_sg4_cmd_attri  [   2:   0]),
  .i8_icb_cmd_beat                (xbar_mg5_ro_to_sg4_cmd_beat   [   1:   0]),
  .i8_icb_cmd_usr                 (xbar_mg5_ro_to_sg4_cmd_usr    [   2:   0]),
  .i8_icb_rsp_ready               (xbar_mg5_ro_to_sg4_rsp_ready             ),
  .i8_icb_rsp_valid               (xbar_mg5_ro_to_sg4_rsp_valid             ),
  .i8_icb_rsp_err                 (xbar_mg5_ro_to_sg4_rsp_err               ),
  .i8_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg4_rsp_excl_ok            ),
  .i8_icb_rsp_rdata               (xbar_mg5_ro_to_sg4_rsp_rdata  [  63:   0]),
  .i8_icb_rsp_usr                 (xbar_mg5_ro_to_sg4_rsp_usr    [   2:   0]),
      .i9_icb_cmd_valid               (xbar_mg5_wo_to_sg4_cmd_valid             ),
  .i9_icb_cmd_ready               (xbar_mg5_wo_to_sg4_cmd_ready             ),
  .i9_icb_cmd_sel                 (xbar_mg5_wo_to_sg4_cmd_sel               ),
  .i9_icb_cmd_read                (xbar_mg5_wo_to_sg4_cmd_read              ),
  .i9_icb_cmd_addr                (xbar_mg5_wo_to_sg4_cmd_addr   [  31:   0]),
  .i9_icb_cmd_wdata               (xbar_mg5_wo_to_sg4_cmd_wdata  [  63:   0]),
  .i9_icb_cmd_wmask               (xbar_mg5_wo_to_sg4_cmd_wmask  [   7:   0]),
  .i9_icb_cmd_size                (xbar_mg5_wo_to_sg4_cmd_size   [   2:   0]),
  .i9_icb_cmd_lock                (xbar_mg5_wo_to_sg4_cmd_lock              ),
  .i9_icb_cmd_excl                (xbar_mg5_wo_to_sg4_cmd_excl              ),
  .i9_icb_cmd_xlen                (xbar_mg5_wo_to_sg4_cmd_xlen   [   7:   0]),
  .i9_icb_cmd_xburst              (xbar_mg5_wo_to_sg4_cmd_xburst [   1:   0]),
  .i9_icb_cmd_modes               (xbar_mg5_wo_to_sg4_cmd_modes  [   1:   0]),
  .i9_icb_cmd_dmode               (xbar_mg5_wo_to_sg4_cmd_dmode             ),
  .i9_icb_cmd_attri               (xbar_mg5_wo_to_sg4_cmd_attri  [   2:   0]),
  .i9_icb_cmd_beat                (xbar_mg5_wo_to_sg4_cmd_beat   [   1:   0]),
  .i9_icb_cmd_usr                 (xbar_mg5_wo_to_sg4_cmd_usr    [   2:   0]),
  .i9_icb_rsp_ready               (xbar_mg5_wo_to_sg4_rsp_ready             ),
  .i9_icb_rsp_valid               (xbar_mg5_wo_to_sg4_rsp_valid             ),
  .i9_icb_rsp_err                 (xbar_mg5_wo_to_sg4_rsp_err               ),
  .i9_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg4_rsp_excl_ok            ),
  .i9_icb_rsp_rdata               (xbar_mg5_wo_to_sg4_rsp_rdata  [  63:   0]),
  .i9_icb_rsp_usr                 (xbar_mg5_wo_to_sg4_rsp_usr    [   2:   0]),
      .i10_icb_cmd_valid              (xbar_mg6_ro_to_sg4_cmd_valid             ),
  .i10_icb_cmd_ready              (xbar_mg6_ro_to_sg4_cmd_ready             ),
  .i10_icb_cmd_sel                (xbar_mg6_ro_to_sg4_cmd_sel               ),
  .i10_icb_cmd_read               (xbar_mg6_ro_to_sg4_cmd_read              ),
  .i10_icb_cmd_addr               (xbar_mg6_ro_to_sg4_cmd_addr   [  31:   0]),
  .i10_icb_cmd_wdata              (xbar_mg6_ro_to_sg4_cmd_wdata  [  63:   0]),
  .i10_icb_cmd_wmask              (xbar_mg6_ro_to_sg4_cmd_wmask  [   7:   0]),
  .i10_icb_cmd_size               (xbar_mg6_ro_to_sg4_cmd_size   [   2:   0]),
  .i10_icb_cmd_lock               (xbar_mg6_ro_to_sg4_cmd_lock              ),
  .i10_icb_cmd_excl               (xbar_mg6_ro_to_sg4_cmd_excl              ),
  .i10_icb_cmd_xlen               (xbar_mg6_ro_to_sg4_cmd_xlen   [   7:   0]),
  .i10_icb_cmd_xburst             (xbar_mg6_ro_to_sg4_cmd_xburst [   1:   0]),
  .i10_icb_cmd_modes              (xbar_mg6_ro_to_sg4_cmd_modes  [   1:   0]),
  .i10_icb_cmd_dmode              (xbar_mg6_ro_to_sg4_cmd_dmode             ),
  .i10_icb_cmd_attri              (xbar_mg6_ro_to_sg4_cmd_attri  [   2:   0]),
  .i10_icb_cmd_beat               (xbar_mg6_ro_to_sg4_cmd_beat   [   1:   0]),
  .i10_icb_cmd_usr                (xbar_mg6_ro_to_sg4_cmd_usr    [   2:   0]),
  .i10_icb_rsp_ready              (xbar_mg6_ro_to_sg4_rsp_ready             ),
  .i10_icb_rsp_valid              (xbar_mg6_ro_to_sg4_rsp_valid             ),
  .i10_icb_rsp_err                (xbar_mg6_ro_to_sg4_rsp_err               ),
  .i10_icb_rsp_excl_ok            (xbar_mg6_ro_to_sg4_rsp_excl_ok            ),
  .i10_icb_rsp_rdata              (xbar_mg6_ro_to_sg4_rsp_rdata  [  63:   0]),
  .i10_icb_rsp_usr                (xbar_mg6_ro_to_sg4_rsp_usr    [   2:   0]),
      .i11_icb_cmd_valid              (xbar_mg6_wo_to_sg4_cmd_valid             ),
  .i11_icb_cmd_ready              (xbar_mg6_wo_to_sg4_cmd_ready             ),
  .i11_icb_cmd_sel                (xbar_mg6_wo_to_sg4_cmd_sel               ),
  .i11_icb_cmd_read               (xbar_mg6_wo_to_sg4_cmd_read              ),
  .i11_icb_cmd_addr               (xbar_mg6_wo_to_sg4_cmd_addr   [  31:   0]),
  .i11_icb_cmd_wdata              (xbar_mg6_wo_to_sg4_cmd_wdata  [  63:   0]),
  .i11_icb_cmd_wmask              (xbar_mg6_wo_to_sg4_cmd_wmask  [   7:   0]),
  .i11_icb_cmd_size               (xbar_mg6_wo_to_sg4_cmd_size   [   2:   0]),
  .i11_icb_cmd_lock               (xbar_mg6_wo_to_sg4_cmd_lock              ),
  .i11_icb_cmd_excl               (xbar_mg6_wo_to_sg4_cmd_excl              ),
  .i11_icb_cmd_xlen               (xbar_mg6_wo_to_sg4_cmd_xlen   [   7:   0]),
  .i11_icb_cmd_xburst             (xbar_mg6_wo_to_sg4_cmd_xburst [   1:   0]),
  .i11_icb_cmd_modes              (xbar_mg6_wo_to_sg4_cmd_modes  [   1:   0]),
  .i11_icb_cmd_dmode              (xbar_mg6_wo_to_sg4_cmd_dmode             ),
  .i11_icb_cmd_attri              (xbar_mg6_wo_to_sg4_cmd_attri  [   2:   0]),
  .i11_icb_cmd_beat               (xbar_mg6_wo_to_sg4_cmd_beat   [   1:   0]),
  .i11_icb_cmd_usr                (xbar_mg6_wo_to_sg4_cmd_usr    [   2:   0]),
  .i11_icb_rsp_ready              (xbar_mg6_wo_to_sg4_rsp_ready             ),
  .i11_icb_rsp_valid              (xbar_mg6_wo_to_sg4_rsp_valid             ),
  .i11_icb_rsp_err                (xbar_mg6_wo_to_sg4_rsp_err               ),
  .i11_icb_rsp_excl_ok            (xbar_mg6_wo_to_sg4_rsp_excl_ok            ),
  .i11_icb_rsp_rdata              (xbar_mg6_wo_to_sg4_rsp_rdata  [  63:   0]),
  .i11_icb_rsp_usr                (xbar_mg6_wo_to_sg4_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
 wire xbar_sg6_rw_arbt_active;
   e603_subsys_xbar_slv6_rw_ficbnto1_bus #(
      .PAYLOAD_NORST(PAYLOAD_NORST),
      .SUPPORT_LOCK(0),
      .I_SUPPORT_RATIO        (0), 
      .O_SUPPORT_RATIO        (0),
      .ICB_FIFO_CMD_DP        (0), 
      .ICB_FIFO_RSP_DP        (0), 
      .ICB_FIFO_CMD_CUT_READY (1),
      .ICB_FIFO_RSP_CUT_READY (1),
      .ARBT_SCHEME         (1),
      .RRBIN_CUT_TIMING       (RRBIN_CUT_TIMING),
      .ARBT_ALLOW_0CYCL_RSP(0),
      .ARBT_FIFO_OUTS_NUM  (8  ),
      .ARBT_FIFO_OUTS_CNT_W(4),
      .ARBT_FIFO_CUT_READY (1) 
   ) u_xbar_sg6_rw_icbnto1(
      .i_clk_en(1'b1),
      .o_clk_en(1'b1),
      .icbnto1_active (xbar_sg6_rw_arbt_active),
      .o_icb_cmd_valid                (slv_grp_6_icb_cmd_valid                  ),
  .o_icb_cmd_ready                (slv_grp_6_icb_cmd_ready                  ),
  .o_icb_cmd_sel                  (slv_grp_6_icb_cmd_sel                    ),
  .o_icb_cmd_read                 (slv_grp_6_icb_cmd_read                   ),
  .o_icb_cmd_addr                 (slv_grp_6_icb_cmd_addr        [  31:   0]),
  .o_icb_cmd_wdata                (slv_grp_6_icb_cmd_wdata       [  63:   0]),
  .o_icb_cmd_wmask                (slv_grp_6_icb_cmd_wmask       [   7:   0]),
  .o_icb_cmd_size                 (slv_grp_6_icb_cmd_size        [   2:   0]),
  .o_icb_cmd_lock                 (slv_grp_6_icb_cmd_lock                   ),
  .o_icb_cmd_excl                 (slv_grp_6_icb_cmd_excl                   ),
  .o_icb_cmd_xlen                 (slv_grp_6_icb_cmd_xlen        [   7:   0]),
  .o_icb_cmd_xburst               (slv_grp_6_icb_cmd_xburst      [   1:   0]),
  .o_icb_cmd_modes                (slv_grp_6_icb_cmd_modes       [   1:   0]),
  .o_icb_cmd_dmode                (slv_grp_6_icb_cmd_dmode                  ),
  .o_icb_cmd_attri                (slv_grp_6_icb_cmd_attri       [   2:   0]),
  .o_icb_cmd_beat                 (slv_grp_6_icb_cmd_beat        [   1:   0]),
  .o_icb_cmd_usr                  (slv_grp_6_icb_cmd_usr         [   2:   0]),
  .o_icb_rsp_ready                (slv_grp_6_icb_rsp_ready                  ),
  .o_icb_rsp_valid                (slv_grp_6_icb_rsp_valid                  ),
  .o_icb_rsp_err                  (slv_grp_6_icb_rsp_err                    ),
  .o_icb_rsp_excl_ok              (slv_grp_6_icb_rsp_excl_ok                ),
  .o_icb_rsp_rdata                (slv_grp_6_icb_rsp_rdata       [  63:   0]),
  .o_icb_rsp_usr                  (slv_grp_6_icb_rsp_usr         [   2:   0]),
      .i0_icb_cmd_valid               (xbar_mg0_ro_to_sg6_cmd_valid             ),
  .i0_icb_cmd_ready               (xbar_mg0_ro_to_sg6_cmd_ready             ),
  .i0_icb_cmd_sel                 (xbar_mg0_ro_to_sg6_cmd_sel               ),
  .i0_icb_cmd_read                (xbar_mg0_ro_to_sg6_cmd_read              ),
  .i0_icb_cmd_addr                (xbar_mg0_ro_to_sg6_cmd_addr   [  31:   0]),
  .i0_icb_cmd_wdata               (xbar_mg0_ro_to_sg6_cmd_wdata  [  63:   0]),
  .i0_icb_cmd_wmask               (xbar_mg0_ro_to_sg6_cmd_wmask  [   7:   0]),
  .i0_icb_cmd_size                (xbar_mg0_ro_to_sg6_cmd_size   [   2:   0]),
  .i0_icb_cmd_lock                (xbar_mg0_ro_to_sg6_cmd_lock              ),
  .i0_icb_cmd_excl                (xbar_mg0_ro_to_sg6_cmd_excl              ),
  .i0_icb_cmd_xlen                (xbar_mg0_ro_to_sg6_cmd_xlen   [   7:   0]),
  .i0_icb_cmd_xburst              (xbar_mg0_ro_to_sg6_cmd_xburst [   1:   0]),
  .i0_icb_cmd_modes               (xbar_mg0_ro_to_sg6_cmd_modes  [   1:   0]),
  .i0_icb_cmd_dmode               (xbar_mg0_ro_to_sg6_cmd_dmode             ),
  .i0_icb_cmd_attri               (xbar_mg0_ro_to_sg6_cmd_attri  [   2:   0]),
  .i0_icb_cmd_beat                (xbar_mg0_ro_to_sg6_cmd_beat   [   1:   0]),
  .i0_icb_cmd_usr                 (xbar_mg0_ro_to_sg6_cmd_usr    [   2:   0]),
  .i0_icb_rsp_ready               (xbar_mg0_ro_to_sg6_rsp_ready             ),
  .i0_icb_rsp_valid               (xbar_mg0_ro_to_sg6_rsp_valid             ),
  .i0_icb_rsp_err                 (xbar_mg0_ro_to_sg6_rsp_err               ),
  .i0_icb_rsp_excl_ok             (xbar_mg0_ro_to_sg6_rsp_excl_ok            ),
  .i0_icb_rsp_rdata               (xbar_mg0_ro_to_sg6_rsp_rdata  [  63:   0]),
  .i0_icb_rsp_usr                 (xbar_mg0_ro_to_sg6_rsp_usr    [   2:   0]),
      .i1_icb_cmd_valid               (xbar_mg0_wo_to_sg6_cmd_valid             ),
  .i1_icb_cmd_ready               (xbar_mg0_wo_to_sg6_cmd_ready             ),
  .i1_icb_cmd_sel                 (xbar_mg0_wo_to_sg6_cmd_sel               ),
  .i1_icb_cmd_read                (xbar_mg0_wo_to_sg6_cmd_read              ),
  .i1_icb_cmd_addr                (xbar_mg0_wo_to_sg6_cmd_addr   [  31:   0]),
  .i1_icb_cmd_wdata               (xbar_mg0_wo_to_sg6_cmd_wdata  [  63:   0]),
  .i1_icb_cmd_wmask               (xbar_mg0_wo_to_sg6_cmd_wmask  [   7:   0]),
  .i1_icb_cmd_size                (xbar_mg0_wo_to_sg6_cmd_size   [   2:   0]),
  .i1_icb_cmd_lock                (xbar_mg0_wo_to_sg6_cmd_lock              ),
  .i1_icb_cmd_excl                (xbar_mg0_wo_to_sg6_cmd_excl              ),
  .i1_icb_cmd_xlen                (xbar_mg0_wo_to_sg6_cmd_xlen   [   7:   0]),
  .i1_icb_cmd_xburst              (xbar_mg0_wo_to_sg6_cmd_xburst [   1:   0]),
  .i1_icb_cmd_modes               (xbar_mg0_wo_to_sg6_cmd_modes  [   1:   0]),
  .i1_icb_cmd_dmode               (xbar_mg0_wo_to_sg6_cmd_dmode             ),
  .i1_icb_cmd_attri               (xbar_mg0_wo_to_sg6_cmd_attri  [   2:   0]),
  .i1_icb_cmd_beat                (xbar_mg0_wo_to_sg6_cmd_beat   [   1:   0]),
  .i1_icb_cmd_usr                 (xbar_mg0_wo_to_sg6_cmd_usr    [   2:   0]),
  .i1_icb_rsp_ready               (xbar_mg0_wo_to_sg6_rsp_ready             ),
  .i1_icb_rsp_valid               (xbar_mg0_wo_to_sg6_rsp_valid             ),
  .i1_icb_rsp_err                 (xbar_mg0_wo_to_sg6_rsp_err               ),
  .i1_icb_rsp_excl_ok             (xbar_mg0_wo_to_sg6_rsp_excl_ok            ),
  .i1_icb_rsp_rdata               (xbar_mg0_wo_to_sg6_rsp_rdata  [  63:   0]),
  .i1_icb_rsp_usr                 (xbar_mg0_wo_to_sg6_rsp_usr    [   2:   0]),
      .i2_icb_cmd_valid               (xbar_mg1_ro_to_sg6_cmd_valid             ),
  .i2_icb_cmd_ready               (xbar_mg1_ro_to_sg6_cmd_ready             ),
  .i2_icb_cmd_sel                 (xbar_mg1_ro_to_sg6_cmd_sel               ),
  .i2_icb_cmd_read                (xbar_mg1_ro_to_sg6_cmd_read              ),
  .i2_icb_cmd_addr                (xbar_mg1_ro_to_sg6_cmd_addr   [  31:   0]),
  .i2_icb_cmd_wdata               (xbar_mg1_ro_to_sg6_cmd_wdata  [  63:   0]),
  .i2_icb_cmd_wmask               (xbar_mg1_ro_to_sg6_cmd_wmask  [   7:   0]),
  .i2_icb_cmd_size                (xbar_mg1_ro_to_sg6_cmd_size   [   2:   0]),
  .i2_icb_cmd_lock                (xbar_mg1_ro_to_sg6_cmd_lock              ),
  .i2_icb_cmd_excl                (xbar_mg1_ro_to_sg6_cmd_excl              ),
  .i2_icb_cmd_xlen                (xbar_mg1_ro_to_sg6_cmd_xlen   [   7:   0]),
  .i2_icb_cmd_xburst              (xbar_mg1_ro_to_sg6_cmd_xburst [   1:   0]),
  .i2_icb_cmd_modes               (xbar_mg1_ro_to_sg6_cmd_modes  [   1:   0]),
  .i2_icb_cmd_dmode               (xbar_mg1_ro_to_sg6_cmd_dmode             ),
  .i2_icb_cmd_attri               (xbar_mg1_ro_to_sg6_cmd_attri  [   2:   0]),
  .i2_icb_cmd_beat                (xbar_mg1_ro_to_sg6_cmd_beat   [   1:   0]),
  .i2_icb_cmd_usr                 (xbar_mg1_ro_to_sg6_cmd_usr    [   2:   0]),
  .i2_icb_rsp_ready               (xbar_mg1_ro_to_sg6_rsp_ready             ),
  .i2_icb_rsp_valid               (xbar_mg1_ro_to_sg6_rsp_valid             ),
  .i2_icb_rsp_err                 (xbar_mg1_ro_to_sg6_rsp_err               ),
  .i2_icb_rsp_excl_ok             (xbar_mg1_ro_to_sg6_rsp_excl_ok            ),
  .i2_icb_rsp_rdata               (xbar_mg1_ro_to_sg6_rsp_rdata  [  63:   0]),
  .i2_icb_rsp_usr                 (xbar_mg1_ro_to_sg6_rsp_usr    [   2:   0]),
      .i3_icb_cmd_valid               (xbar_mg2_wo_to_sg6_cmd_valid             ),
  .i3_icb_cmd_ready               (xbar_mg2_wo_to_sg6_cmd_ready             ),
  .i3_icb_cmd_sel                 (xbar_mg2_wo_to_sg6_cmd_sel               ),
  .i3_icb_cmd_read                (xbar_mg2_wo_to_sg6_cmd_read              ),
  .i3_icb_cmd_addr                (xbar_mg2_wo_to_sg6_cmd_addr   [  31:   0]),
  .i3_icb_cmd_wdata               (xbar_mg2_wo_to_sg6_cmd_wdata  [  63:   0]),
  .i3_icb_cmd_wmask               (xbar_mg2_wo_to_sg6_cmd_wmask  [   7:   0]),
  .i3_icb_cmd_size                (xbar_mg2_wo_to_sg6_cmd_size   [   2:   0]),
  .i3_icb_cmd_lock                (xbar_mg2_wo_to_sg6_cmd_lock              ),
  .i3_icb_cmd_excl                (xbar_mg2_wo_to_sg6_cmd_excl              ),
  .i3_icb_cmd_xlen                (xbar_mg2_wo_to_sg6_cmd_xlen   [   7:   0]),
  .i3_icb_cmd_xburst              (xbar_mg2_wo_to_sg6_cmd_xburst [   1:   0]),
  .i3_icb_cmd_modes               (xbar_mg2_wo_to_sg6_cmd_modes  [   1:   0]),
  .i3_icb_cmd_dmode               (xbar_mg2_wo_to_sg6_cmd_dmode             ),
  .i3_icb_cmd_attri               (xbar_mg2_wo_to_sg6_cmd_attri  [   2:   0]),
  .i3_icb_cmd_beat                (xbar_mg2_wo_to_sg6_cmd_beat   [   1:   0]),
  .i3_icb_cmd_usr                 (xbar_mg2_wo_to_sg6_cmd_usr    [   2:   0]),
  .i3_icb_rsp_ready               (xbar_mg2_wo_to_sg6_rsp_ready             ),
  .i3_icb_rsp_valid               (xbar_mg2_wo_to_sg6_rsp_valid             ),
  .i3_icb_rsp_err                 (xbar_mg2_wo_to_sg6_rsp_err               ),
  .i3_icb_rsp_excl_ok             (xbar_mg2_wo_to_sg6_rsp_excl_ok            ),
  .i3_icb_rsp_rdata               (xbar_mg2_wo_to_sg6_rsp_rdata  [  63:   0]),
  .i3_icb_rsp_usr                 (xbar_mg2_wo_to_sg6_rsp_usr    [   2:   0]),
      .i4_icb_cmd_valid               (xbar_mg3_ro_to_sg6_cmd_valid             ),
  .i4_icb_cmd_ready               (xbar_mg3_ro_to_sg6_cmd_ready             ),
  .i4_icb_cmd_sel                 (xbar_mg3_ro_to_sg6_cmd_sel               ),
  .i4_icb_cmd_read                (xbar_mg3_ro_to_sg6_cmd_read              ),
  .i4_icb_cmd_addr                (xbar_mg3_ro_to_sg6_cmd_addr   [  31:   0]),
  .i4_icb_cmd_wdata               (xbar_mg3_ro_to_sg6_cmd_wdata  [  63:   0]),
  .i4_icb_cmd_wmask               (xbar_mg3_ro_to_sg6_cmd_wmask  [   7:   0]),
  .i4_icb_cmd_size                (xbar_mg3_ro_to_sg6_cmd_size   [   2:   0]),
  .i4_icb_cmd_lock                (xbar_mg3_ro_to_sg6_cmd_lock              ),
  .i4_icb_cmd_excl                (xbar_mg3_ro_to_sg6_cmd_excl              ),
  .i4_icb_cmd_xlen                (xbar_mg3_ro_to_sg6_cmd_xlen   [   7:   0]),
  .i4_icb_cmd_xburst              (xbar_mg3_ro_to_sg6_cmd_xburst [   1:   0]),
  .i4_icb_cmd_modes               (xbar_mg3_ro_to_sg6_cmd_modes  [   1:   0]),
  .i4_icb_cmd_dmode               (xbar_mg3_ro_to_sg6_cmd_dmode             ),
  .i4_icb_cmd_attri               (xbar_mg3_ro_to_sg6_cmd_attri  [   2:   0]),
  .i4_icb_cmd_beat                (xbar_mg3_ro_to_sg6_cmd_beat   [   1:   0]),
  .i4_icb_cmd_usr                 (xbar_mg3_ro_to_sg6_cmd_usr    [   2:   0]),
  .i4_icb_rsp_ready               (xbar_mg3_ro_to_sg6_rsp_ready             ),
  .i4_icb_rsp_valid               (xbar_mg3_ro_to_sg6_rsp_valid             ),
  .i4_icb_rsp_err                 (xbar_mg3_ro_to_sg6_rsp_err               ),
  .i4_icb_rsp_excl_ok             (xbar_mg3_ro_to_sg6_rsp_excl_ok            ),
  .i4_icb_rsp_rdata               (xbar_mg3_ro_to_sg6_rsp_rdata  [  63:   0]),
  .i4_icb_rsp_usr                 (xbar_mg3_ro_to_sg6_rsp_usr    [   2:   0]),
      .i5_icb_cmd_valid               (xbar_mg3_wo_to_sg6_cmd_valid             ),
  .i5_icb_cmd_ready               (xbar_mg3_wo_to_sg6_cmd_ready             ),
  .i5_icb_cmd_sel                 (xbar_mg3_wo_to_sg6_cmd_sel               ),
  .i5_icb_cmd_read                (xbar_mg3_wo_to_sg6_cmd_read              ),
  .i5_icb_cmd_addr                (xbar_mg3_wo_to_sg6_cmd_addr   [  31:   0]),
  .i5_icb_cmd_wdata               (xbar_mg3_wo_to_sg6_cmd_wdata  [  63:   0]),
  .i5_icb_cmd_wmask               (xbar_mg3_wo_to_sg6_cmd_wmask  [   7:   0]),
  .i5_icb_cmd_size                (xbar_mg3_wo_to_sg6_cmd_size   [   2:   0]),
  .i5_icb_cmd_lock                (xbar_mg3_wo_to_sg6_cmd_lock              ),
  .i5_icb_cmd_excl                (xbar_mg3_wo_to_sg6_cmd_excl              ),
  .i5_icb_cmd_xlen                (xbar_mg3_wo_to_sg6_cmd_xlen   [   7:   0]),
  .i5_icb_cmd_xburst              (xbar_mg3_wo_to_sg6_cmd_xburst [   1:   0]),
  .i5_icb_cmd_modes               (xbar_mg3_wo_to_sg6_cmd_modes  [   1:   0]),
  .i5_icb_cmd_dmode               (xbar_mg3_wo_to_sg6_cmd_dmode             ),
  .i5_icb_cmd_attri               (xbar_mg3_wo_to_sg6_cmd_attri  [   2:   0]),
  .i5_icb_cmd_beat                (xbar_mg3_wo_to_sg6_cmd_beat   [   1:   0]),
  .i5_icb_cmd_usr                 (xbar_mg3_wo_to_sg6_cmd_usr    [   2:   0]),
  .i5_icb_rsp_ready               (xbar_mg3_wo_to_sg6_rsp_ready             ),
  .i5_icb_rsp_valid               (xbar_mg3_wo_to_sg6_rsp_valid             ),
  .i5_icb_rsp_err                 (xbar_mg3_wo_to_sg6_rsp_err               ),
  .i5_icb_rsp_excl_ok             (xbar_mg3_wo_to_sg6_rsp_excl_ok            ),
  .i5_icb_rsp_rdata               (xbar_mg3_wo_to_sg6_rsp_rdata  [  63:   0]),
  .i5_icb_rsp_usr                 (xbar_mg3_wo_to_sg6_rsp_usr    [   2:   0]),
      .i6_icb_cmd_valid               (xbar_mg4_ro_to_sg6_cmd_valid             ),
  .i6_icb_cmd_ready               (xbar_mg4_ro_to_sg6_cmd_ready             ),
  .i6_icb_cmd_sel                 (xbar_mg4_ro_to_sg6_cmd_sel               ),
  .i6_icb_cmd_read                (xbar_mg4_ro_to_sg6_cmd_read              ),
  .i6_icb_cmd_addr                (xbar_mg4_ro_to_sg6_cmd_addr   [  31:   0]),
  .i6_icb_cmd_wdata               (xbar_mg4_ro_to_sg6_cmd_wdata  [  63:   0]),
  .i6_icb_cmd_wmask               (xbar_mg4_ro_to_sg6_cmd_wmask  [   7:   0]),
  .i6_icb_cmd_size                (xbar_mg4_ro_to_sg6_cmd_size   [   2:   0]),
  .i6_icb_cmd_lock                (xbar_mg4_ro_to_sg6_cmd_lock              ),
  .i6_icb_cmd_excl                (xbar_mg4_ro_to_sg6_cmd_excl              ),
  .i6_icb_cmd_xlen                (xbar_mg4_ro_to_sg6_cmd_xlen   [   7:   0]),
  .i6_icb_cmd_xburst              (xbar_mg4_ro_to_sg6_cmd_xburst [   1:   0]),
  .i6_icb_cmd_modes               (xbar_mg4_ro_to_sg6_cmd_modes  [   1:   0]),
  .i6_icb_cmd_dmode               (xbar_mg4_ro_to_sg6_cmd_dmode             ),
  .i6_icb_cmd_attri               (xbar_mg4_ro_to_sg6_cmd_attri  [   2:   0]),
  .i6_icb_cmd_beat                (xbar_mg4_ro_to_sg6_cmd_beat   [   1:   0]),
  .i6_icb_cmd_usr                 (xbar_mg4_ro_to_sg6_cmd_usr    [   2:   0]),
  .i6_icb_rsp_ready               (xbar_mg4_ro_to_sg6_rsp_ready             ),
  .i6_icb_rsp_valid               (xbar_mg4_ro_to_sg6_rsp_valid             ),
  .i6_icb_rsp_err                 (xbar_mg4_ro_to_sg6_rsp_err               ),
  .i6_icb_rsp_excl_ok             (xbar_mg4_ro_to_sg6_rsp_excl_ok            ),
  .i6_icb_rsp_rdata               (xbar_mg4_ro_to_sg6_rsp_rdata  [  63:   0]),
  .i6_icb_rsp_usr                 (xbar_mg4_ro_to_sg6_rsp_usr    [   2:   0]),
      .i7_icb_cmd_valid               (xbar_mg4_wo_to_sg6_cmd_valid             ),
  .i7_icb_cmd_ready               (xbar_mg4_wo_to_sg6_cmd_ready             ),
  .i7_icb_cmd_sel                 (xbar_mg4_wo_to_sg6_cmd_sel               ),
  .i7_icb_cmd_read                (xbar_mg4_wo_to_sg6_cmd_read              ),
  .i7_icb_cmd_addr                (xbar_mg4_wo_to_sg6_cmd_addr   [  31:   0]),
  .i7_icb_cmd_wdata               (xbar_mg4_wo_to_sg6_cmd_wdata  [  63:   0]),
  .i7_icb_cmd_wmask               (xbar_mg4_wo_to_sg6_cmd_wmask  [   7:   0]),
  .i7_icb_cmd_size                (xbar_mg4_wo_to_sg6_cmd_size   [   2:   0]),
  .i7_icb_cmd_lock                (xbar_mg4_wo_to_sg6_cmd_lock              ),
  .i7_icb_cmd_excl                (xbar_mg4_wo_to_sg6_cmd_excl              ),
  .i7_icb_cmd_xlen                (xbar_mg4_wo_to_sg6_cmd_xlen   [   7:   0]),
  .i7_icb_cmd_xburst              (xbar_mg4_wo_to_sg6_cmd_xburst [   1:   0]),
  .i7_icb_cmd_modes               (xbar_mg4_wo_to_sg6_cmd_modes  [   1:   0]),
  .i7_icb_cmd_dmode               (xbar_mg4_wo_to_sg6_cmd_dmode             ),
  .i7_icb_cmd_attri               (xbar_mg4_wo_to_sg6_cmd_attri  [   2:   0]),
  .i7_icb_cmd_beat                (xbar_mg4_wo_to_sg6_cmd_beat   [   1:   0]),
  .i7_icb_cmd_usr                 (xbar_mg4_wo_to_sg6_cmd_usr    [   2:   0]),
  .i7_icb_rsp_ready               (xbar_mg4_wo_to_sg6_rsp_ready             ),
  .i7_icb_rsp_valid               (xbar_mg4_wo_to_sg6_rsp_valid             ),
  .i7_icb_rsp_err                 (xbar_mg4_wo_to_sg6_rsp_err               ),
  .i7_icb_rsp_excl_ok             (xbar_mg4_wo_to_sg6_rsp_excl_ok            ),
  .i7_icb_rsp_rdata               (xbar_mg4_wo_to_sg6_rsp_rdata  [  63:   0]),
  .i7_icb_rsp_usr                 (xbar_mg4_wo_to_sg6_rsp_usr    [   2:   0]),
      .i8_icb_cmd_valid               (xbar_mg5_ro_to_sg6_cmd_valid             ),
  .i8_icb_cmd_ready               (xbar_mg5_ro_to_sg6_cmd_ready             ),
  .i8_icb_cmd_sel                 (xbar_mg5_ro_to_sg6_cmd_sel               ),
  .i8_icb_cmd_read                (xbar_mg5_ro_to_sg6_cmd_read              ),
  .i8_icb_cmd_addr                (xbar_mg5_ro_to_sg6_cmd_addr   [  31:   0]),
  .i8_icb_cmd_wdata               (xbar_mg5_ro_to_sg6_cmd_wdata  [  63:   0]),
  .i8_icb_cmd_wmask               (xbar_mg5_ro_to_sg6_cmd_wmask  [   7:   0]),
  .i8_icb_cmd_size                (xbar_mg5_ro_to_sg6_cmd_size   [   2:   0]),
  .i8_icb_cmd_lock                (xbar_mg5_ro_to_sg6_cmd_lock              ),
  .i8_icb_cmd_excl                (xbar_mg5_ro_to_sg6_cmd_excl              ),
  .i8_icb_cmd_xlen                (xbar_mg5_ro_to_sg6_cmd_xlen   [   7:   0]),
  .i8_icb_cmd_xburst              (xbar_mg5_ro_to_sg6_cmd_xburst [   1:   0]),
  .i8_icb_cmd_modes               (xbar_mg5_ro_to_sg6_cmd_modes  [   1:   0]),
  .i8_icb_cmd_dmode               (xbar_mg5_ro_to_sg6_cmd_dmode             ),
  .i8_icb_cmd_attri               (xbar_mg5_ro_to_sg6_cmd_attri  [   2:   0]),
  .i8_icb_cmd_beat                (xbar_mg5_ro_to_sg6_cmd_beat   [   1:   0]),
  .i8_icb_cmd_usr                 (xbar_mg5_ro_to_sg6_cmd_usr    [   2:   0]),
  .i8_icb_rsp_ready               (xbar_mg5_ro_to_sg6_rsp_ready             ),
  .i8_icb_rsp_valid               (xbar_mg5_ro_to_sg6_rsp_valid             ),
  .i8_icb_rsp_err                 (xbar_mg5_ro_to_sg6_rsp_err               ),
  .i8_icb_rsp_excl_ok             (xbar_mg5_ro_to_sg6_rsp_excl_ok            ),
  .i8_icb_rsp_rdata               (xbar_mg5_ro_to_sg6_rsp_rdata  [  63:   0]),
  .i8_icb_rsp_usr                 (xbar_mg5_ro_to_sg6_rsp_usr    [   2:   0]),
      .i9_icb_cmd_valid               (xbar_mg5_wo_to_sg6_cmd_valid             ),
  .i9_icb_cmd_ready               (xbar_mg5_wo_to_sg6_cmd_ready             ),
  .i9_icb_cmd_sel                 (xbar_mg5_wo_to_sg6_cmd_sel               ),
  .i9_icb_cmd_read                (xbar_mg5_wo_to_sg6_cmd_read              ),
  .i9_icb_cmd_addr                (xbar_mg5_wo_to_sg6_cmd_addr   [  31:   0]),
  .i9_icb_cmd_wdata               (xbar_mg5_wo_to_sg6_cmd_wdata  [  63:   0]),
  .i9_icb_cmd_wmask               (xbar_mg5_wo_to_sg6_cmd_wmask  [   7:   0]),
  .i9_icb_cmd_size                (xbar_mg5_wo_to_sg6_cmd_size   [   2:   0]),
  .i9_icb_cmd_lock                (xbar_mg5_wo_to_sg6_cmd_lock              ),
  .i9_icb_cmd_excl                (xbar_mg5_wo_to_sg6_cmd_excl              ),
  .i9_icb_cmd_xlen                (xbar_mg5_wo_to_sg6_cmd_xlen   [   7:   0]),
  .i9_icb_cmd_xburst              (xbar_mg5_wo_to_sg6_cmd_xburst [   1:   0]),
  .i9_icb_cmd_modes               (xbar_mg5_wo_to_sg6_cmd_modes  [   1:   0]),
  .i9_icb_cmd_dmode               (xbar_mg5_wo_to_sg6_cmd_dmode             ),
  .i9_icb_cmd_attri               (xbar_mg5_wo_to_sg6_cmd_attri  [   2:   0]),
  .i9_icb_cmd_beat                (xbar_mg5_wo_to_sg6_cmd_beat   [   1:   0]),
  .i9_icb_cmd_usr                 (xbar_mg5_wo_to_sg6_cmd_usr    [   2:   0]),
  .i9_icb_rsp_ready               (xbar_mg5_wo_to_sg6_rsp_ready             ),
  .i9_icb_rsp_valid               (xbar_mg5_wo_to_sg6_rsp_valid             ),
  .i9_icb_rsp_err                 (xbar_mg5_wo_to_sg6_rsp_err               ),
  .i9_icb_rsp_excl_ok             (xbar_mg5_wo_to_sg6_rsp_excl_ok            ),
  .i9_icb_rsp_rdata               (xbar_mg5_wo_to_sg6_rsp_rdata  [  63:   0]),
  .i9_icb_rsp_usr                 (xbar_mg5_wo_to_sg6_rsp_usr    [   2:   0]),
      .i10_icb_cmd_valid              (xbar_mg6_ro_to_sg6_cmd_valid             ),
  .i10_icb_cmd_ready              (xbar_mg6_ro_to_sg6_cmd_ready             ),
  .i10_icb_cmd_sel                (xbar_mg6_ro_to_sg6_cmd_sel               ),
  .i10_icb_cmd_read               (xbar_mg6_ro_to_sg6_cmd_read              ),
  .i10_icb_cmd_addr               (xbar_mg6_ro_to_sg6_cmd_addr   [  31:   0]),
  .i10_icb_cmd_wdata              (xbar_mg6_ro_to_sg6_cmd_wdata  [  63:   0]),
  .i10_icb_cmd_wmask              (xbar_mg6_ro_to_sg6_cmd_wmask  [   7:   0]),
  .i10_icb_cmd_size               (xbar_mg6_ro_to_sg6_cmd_size   [   2:   0]),
  .i10_icb_cmd_lock               (xbar_mg6_ro_to_sg6_cmd_lock              ),
  .i10_icb_cmd_excl               (xbar_mg6_ro_to_sg6_cmd_excl              ),
  .i10_icb_cmd_xlen               (xbar_mg6_ro_to_sg6_cmd_xlen   [   7:   0]),
  .i10_icb_cmd_xburst             (xbar_mg6_ro_to_sg6_cmd_xburst [   1:   0]),
  .i10_icb_cmd_modes              (xbar_mg6_ro_to_sg6_cmd_modes  [   1:   0]),
  .i10_icb_cmd_dmode              (xbar_mg6_ro_to_sg6_cmd_dmode             ),
  .i10_icb_cmd_attri              (xbar_mg6_ro_to_sg6_cmd_attri  [   2:   0]),
  .i10_icb_cmd_beat               (xbar_mg6_ro_to_sg6_cmd_beat   [   1:   0]),
  .i10_icb_cmd_usr                (xbar_mg6_ro_to_sg6_cmd_usr    [   2:   0]),
  .i10_icb_rsp_ready              (xbar_mg6_ro_to_sg6_rsp_ready             ),
  .i10_icb_rsp_valid              (xbar_mg6_ro_to_sg6_rsp_valid             ),
  .i10_icb_rsp_err                (xbar_mg6_ro_to_sg6_rsp_err               ),
  .i10_icb_rsp_excl_ok            (xbar_mg6_ro_to_sg6_rsp_excl_ok            ),
  .i10_icb_rsp_rdata              (xbar_mg6_ro_to_sg6_rsp_rdata  [  63:   0]),
  .i10_icb_rsp_usr                (xbar_mg6_ro_to_sg6_rsp_usr    [   2:   0]),
      .i11_icb_cmd_valid              (xbar_mg6_wo_to_sg6_cmd_valid             ),
  .i11_icb_cmd_ready              (xbar_mg6_wo_to_sg6_cmd_ready             ),
  .i11_icb_cmd_sel                (xbar_mg6_wo_to_sg6_cmd_sel               ),
  .i11_icb_cmd_read               (xbar_mg6_wo_to_sg6_cmd_read              ),
  .i11_icb_cmd_addr               (xbar_mg6_wo_to_sg6_cmd_addr   [  31:   0]),
  .i11_icb_cmd_wdata              (xbar_mg6_wo_to_sg6_cmd_wdata  [  63:   0]),
  .i11_icb_cmd_wmask              (xbar_mg6_wo_to_sg6_cmd_wmask  [   7:   0]),
  .i11_icb_cmd_size               (xbar_mg6_wo_to_sg6_cmd_size   [   2:   0]),
  .i11_icb_cmd_lock               (xbar_mg6_wo_to_sg6_cmd_lock              ),
  .i11_icb_cmd_excl               (xbar_mg6_wo_to_sg6_cmd_excl              ),
  .i11_icb_cmd_xlen               (xbar_mg6_wo_to_sg6_cmd_xlen   [   7:   0]),
  .i11_icb_cmd_xburst             (xbar_mg6_wo_to_sg6_cmd_xburst [   1:   0]),
  .i11_icb_cmd_modes              (xbar_mg6_wo_to_sg6_cmd_modes  [   1:   0]),
  .i11_icb_cmd_dmode              (xbar_mg6_wo_to_sg6_cmd_dmode             ),
  .i11_icb_cmd_attri              (xbar_mg6_wo_to_sg6_cmd_attri  [   2:   0]),
  .i11_icb_cmd_beat               (xbar_mg6_wo_to_sg6_cmd_beat   [   1:   0]),
  .i11_icb_cmd_usr                (xbar_mg6_wo_to_sg6_cmd_usr    [   2:   0]),
  .i11_icb_rsp_ready              (xbar_mg6_wo_to_sg6_rsp_ready             ),
  .i11_icb_rsp_valid              (xbar_mg6_wo_to_sg6_rsp_valid             ),
  .i11_icb_rsp_err                (xbar_mg6_wo_to_sg6_rsp_err               ),
  .i11_icb_rsp_excl_ok            (xbar_mg6_wo_to_sg6_rsp_excl_ok            ),
  .i11_icb_rsp_rdata              (xbar_mg6_wo_to_sg6_rsp_rdata  [  63:   0]),
  .i11_icb_rsp_usr                (xbar_mg6_wo_to_sg6_rsp_usr    [   2:   0]),
    .clk  (clk_fab  ),
    .rst_n(rst_n)
  );
  wire fab_active_pre = 1'b0
         | i_axi_bus_active 
         | udma_r_icb_bus_active 
         | udma_w_icb_bus_active 
         | dummy_icb_bus_active 
         | dummy_axi_bus_active 
         | dummy_ahbl_bus_active 
         | eth_axi_bus_active 
         | biu2iram_icb_bus_pend_active
         | biu2dram_icb_bus_pend_active
         | addr0_icb_bus_pend_active
         | qspi0_ro_icb_bus_pend_active
         | eth_cfg_apb_bus_pend_active
         | biu2ppi_icb_bus_pend_active
         | o0_axi_bus_pend_active
         | dummy_slv_icb_bus_pend_active
   ;
  wire fab_icb_any_active = 1'b0
         | i_axi_bus_active 
         | udma_r_icb_bus_active 
         | udma_w_icb_bus_active 
         | dummy_icb_bus_active 
         | dummy_axi_bus_active 
         | dummy_ahbl_bus_active 
         | eth_axi_bus_active 
         | biu2iram_icb_bus_icb_active
         | biu2dram_icb_bus_icb_active
         | addr0_icb_bus_icb_active
         | qspi0_ro_icb_bus_icb_active
         | eth_cfg_apb_bus_icb_active
         | biu2ppi_icb_bus_icb_active
         | o0_axi_bus_icb_active
         | dummy_slv_icb_bus_icb_active
   ;
     wire fab_active_d1_r; 
     wire fab_active_d2_r;
     wire fab_active_d3_r;
     wire fab_active_d4_r;
     wire fab_active_d1_nxt = fab_active_pre; 
     wire fab_active_d2_nxt = fab_active_d1_r;
     wire fab_active_d3_nxt = fab_active_d2_r;
     wire fab_active_d4_nxt = fab_active_d3_r;
     wire fab_active_d1_ena = (fab_active_d1_nxt ^ fab_active_d1_r);
e603_gnrl_dfflr #(1) fab_active_d1_dfflr (fab_active_d1_ena, fab_active_d1_nxt, fab_active_d1_r, clk, rst_n);// VPP_NO_REG_PARSE
     wire fab_active_d2_ena = (fab_active_d2_nxt ^ fab_active_d2_r);
e603_gnrl_dfflr #(1) fab_active_d2_dfflr (fab_active_d2_ena, fab_active_d2_nxt, fab_active_d2_r, clk, rst_n);// VPP_NO_REG_PARSE
     wire fab_active_d3_ena = (fab_active_d3_nxt ^ fab_active_d3_r);
e603_gnrl_dfflr #(1) fab_active_d3_dfflr (fab_active_d3_ena, fab_active_d3_nxt, fab_active_d3_r, clk, rst_n);// VPP_NO_REG_PARSE
     wire fab_active_d4_ena = (fab_active_d4_nxt ^ fab_active_d4_r);
e603_gnrl_dfflr #(1) fab_active_d4_dfflr (fab_active_d4_ena, fab_active_d4_nxt, fab_active_d4_r, clk, rst_n);// VPP_NO_REG_PARSE
    assign fab_active = fab_active_pre 
                      | fab_active_d1_r 
                      | fab_active_d2_r
                      | fab_active_d3_r
                      | fab_active_d4_r
                      ;
endmodule
module e603_subsys_xbar_mst0_ro_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
        .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata({(64){1'b0}}),
    .i_icb_cmd_wmask({(64/8){1'b0}}),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 447:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst1_ro_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
        .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata({(64){1'b0}}),
    .i_icb_cmd_wmask({(64/8){1'b0}}),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 447:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst2_ro_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
        .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata({(64){1'b0}}),
    .i_icb_cmd_wmask({(64/8){1'b0}}),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 447:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst3_ro_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
        .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata({(64){1'b0}}),
    .i_icb_cmd_wmask({(64/8){1'b0}}),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 447:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst4_ro_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
        .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata({(64){1'b0}}),
    .i_icb_cmd_wmask({(64/8){1'b0}}),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 447:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst5_ro_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
        .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata({(64){1'b0}}),
    .i_icb_cmd_wmask({(64/8){1'b0}}),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 447:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst6_ro_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
        .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata({(64){1'b0}}),
    .i_icb_cmd_wmask({(64/8){1'b0}}),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 447:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst0_wo_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .o_bus_icb_rsp_rdata({(64*7){1'b0}}),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst1_wo_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .o_bus_icb_rsp_rdata({(64*7){1'b0}}),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst2_wo_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .o_bus_icb_rsp_rdata({(64*7){1'b0}}),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst3_wo_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .o_bus_icb_rsp_rdata({(64*7){1'b0}}),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst4_wo_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .o_bus_icb_rsp_rdata({(64*7){1'b0}}),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst5_wo_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .o_bus_icb_rsp_rdata({(64*7){1'b0}}),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_mst6_wo_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter O3_BASE_ADDR       = 32'h0,       
  parameter O3_BASE_REGION_LSB = 12,
  parameter O4_BASE_ADDR       = 32'h0,       
  parameter O4_BASE_REGION_LSB = 12,
  parameter O5_BASE_ADDR       = 32'h0,       
  parameter O5_BASE_REGION_LSB = 12,
  parameter O6_BASE_ADDR       = 32'h0,       
  parameter O6_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input                          o2_icb_enable,
    output             o2_icb_cmd_valid              ,
  input              o2_icb_cmd_ready              ,
  output             o2_icb_cmd_sel                ,
  output             o2_icb_cmd_read               ,
  output [  31:   0] o2_icb_cmd_addr               ,
  output [  63:   0] o2_icb_cmd_wdata              ,
  output [   7:   0] o2_icb_cmd_wmask              ,
  output [   2:   0] o2_icb_cmd_size               ,
  output             o2_icb_cmd_lock               ,
  output             o2_icb_cmd_excl               ,
  output [   7:   0] o2_icb_cmd_xlen               ,
  output [   1:   0] o2_icb_cmd_xburst             ,
  output [   1:   0] o2_icb_cmd_modes              ,
  output             o2_icb_cmd_dmode              ,
  output [   2:   0] o2_icb_cmd_attri              ,
  output [   1:   0] o2_icb_cmd_beat               ,
  output [   2:   0] o2_icb_cmd_usr                ,
  output             o2_icb_rsp_ready              ,
  input              o2_icb_rsp_valid              ,
  input              o2_icb_rsp_err                ,
  input              o2_icb_rsp_excl_ok            ,
  input  [  63:   0] o2_icb_rsp_rdata              ,
  input  [   2:   0] o2_icb_rsp_usr                ,
  input                          o3_icb_enable,
    output             o3_icb_cmd_valid              ,
  input              o3_icb_cmd_ready              ,
  output             o3_icb_cmd_sel                ,
  output             o3_icb_cmd_read               ,
  output [  31:   0] o3_icb_cmd_addr               ,
  output [  63:   0] o3_icb_cmd_wdata              ,
  output [   7:   0] o3_icb_cmd_wmask              ,
  output [   2:   0] o3_icb_cmd_size               ,
  output             o3_icb_cmd_lock               ,
  output             o3_icb_cmd_excl               ,
  output [   7:   0] o3_icb_cmd_xlen               ,
  output [   1:   0] o3_icb_cmd_xburst             ,
  output [   1:   0] o3_icb_cmd_modes              ,
  output             o3_icb_cmd_dmode              ,
  output [   2:   0] o3_icb_cmd_attri              ,
  output [   1:   0] o3_icb_cmd_beat               ,
  output [   2:   0] o3_icb_cmd_usr                ,
  output             o3_icb_rsp_ready              ,
  input              o3_icb_rsp_valid              ,
  input              o3_icb_rsp_err                ,
  input              o3_icb_rsp_excl_ok            ,
  input  [  63:   0] o3_icb_rsp_rdata              ,
  input  [   2:   0] o3_icb_rsp_usr                ,
  input                          o4_icb_enable,
    output             o4_icb_cmd_valid              ,
  input              o4_icb_cmd_ready              ,
  output             o4_icb_cmd_sel                ,
  output             o4_icb_cmd_read               ,
  output [  31:   0] o4_icb_cmd_addr               ,
  output [  63:   0] o4_icb_cmd_wdata              ,
  output [   7:   0] o4_icb_cmd_wmask              ,
  output [   2:   0] o4_icb_cmd_size               ,
  output             o4_icb_cmd_lock               ,
  output             o4_icb_cmd_excl               ,
  output [   7:   0] o4_icb_cmd_xlen               ,
  output [   1:   0] o4_icb_cmd_xburst             ,
  output [   1:   0] o4_icb_cmd_modes              ,
  output             o4_icb_cmd_dmode              ,
  output [   2:   0] o4_icb_cmd_attri              ,
  output [   1:   0] o4_icb_cmd_beat               ,
  output [   2:   0] o4_icb_cmd_usr                ,
  output             o4_icb_rsp_ready              ,
  input              o4_icb_rsp_valid              ,
  input              o4_icb_rsp_err                ,
  input              o4_icb_rsp_excl_ok            ,
  input  [  63:   0] o4_icb_rsp_rdata              ,
  input  [   2:   0] o4_icb_rsp_usr                ,
  input                          o5_icb_enable,
    output             o5_icb_cmd_valid              ,
  input              o5_icb_cmd_ready              ,
  output             o5_icb_cmd_sel                ,
  output             o5_icb_cmd_read               ,
  output [  31:   0] o5_icb_cmd_addr               ,
  output [  63:   0] o5_icb_cmd_wdata              ,
  output [   7:   0] o5_icb_cmd_wmask              ,
  output [   2:   0] o5_icb_cmd_size               ,
  output             o5_icb_cmd_lock               ,
  output             o5_icb_cmd_excl               ,
  output [   7:   0] o5_icb_cmd_xlen               ,
  output [   1:   0] o5_icb_cmd_xburst             ,
  output [   1:   0] o5_icb_cmd_modes              ,
  output             o5_icb_cmd_dmode              ,
  output [   2:   0] o5_icb_cmd_attri              ,
  output [   1:   0] o5_icb_cmd_beat               ,
  output [   2:   0] o5_icb_cmd_usr                ,
  output             o5_icb_rsp_ready              ,
  input              o5_icb_rsp_valid              ,
  input              o5_icb_rsp_err                ,
  input              o5_icb_rsp_excl_ok            ,
  input  [  63:   0] o5_icb_rsp_rdata              ,
  input  [   2:   0] o5_icb_rsp_usr                ,
    output             o6_icb_cmd_valid              ,
  input              o6_icb_cmd_ready              ,
  output             o6_icb_cmd_sel                ,
  output             o6_icb_cmd_read               ,
  output [  31:   0] o6_icb_cmd_addr               ,
  output [  63:   0] o6_icb_cmd_wdata              ,
  output [   7:   0] o6_icb_cmd_wmask              ,
  output [   2:   0] o6_icb_cmd_size               ,
  output             o6_icb_cmd_lock               ,
  output             o6_icb_cmd_excl               ,
  output [   7:   0] o6_icb_cmd_xlen               ,
  output [   1:   0] o6_icb_cmd_xburst             ,
  output [   1:   0] o6_icb_cmd_modes              ,
  output             o6_icb_cmd_dmode              ,
  output [   2:   0] o6_icb_cmd_attri              ,
  output [   1:   0] o6_icb_cmd_beat               ,
  output [   2:   0] o6_icb_cmd_usr                ,
  output             o6_icb_rsp_ready              ,
  input              o6_icb_rsp_valid              ,
  input              o6_icb_rsp_err                ,
  input              o6_icb_rsp_excl_ok            ,
  input  [  63:   0] o6_icb_rsp_rdata              ,
  input  [   2:   0] o6_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   6:   0] splt_bus_icb_cmd_valid        ;
  wire    [   6:   0] splt_bus_icb_cmd_ready        ;
  wire    [   6:   0] splt_bus_icb_cmd_sel          ;
  wire    [   6:   0] splt_bus_icb_cmd_read         ;
  wire    [ 223:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 447:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  55:   0] splt_bus_icb_cmd_wmask        ;
  wire    [  20:   0] splt_bus_icb_cmd_size         ;
  wire    [   6:   0] splt_bus_icb_cmd_lock         ;
  wire    [   6:   0] splt_bus_icb_cmd_excl         ;
  wire    [  55:   0] splt_bus_icb_cmd_xlen         ;
  wire    [  13:   0] splt_bus_icb_cmd_xburst       ;
  wire    [  13:   0] splt_bus_icb_cmd_modes        ;
  wire    [   6:   0] splt_bus_icb_cmd_dmode        ;
  wire    [  20:   0] splt_bus_icb_cmd_attri        ;
  wire    [  13:   0] splt_bus_icb_cmd_beat         ;
  wire    [  20:   0] splt_bus_icb_cmd_usr          ;
  wire    [   6:   0] splt_bus_icb_rsp_ready        ;
  wire    [   6:   0] splt_bus_icb_rsp_valid        ;
  wire    [   6:   0] splt_bus_icb_rsp_err          ;
  wire    [   6:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 447:   0] splt_bus_icb_rsp_rdata        ;
  wire    [  20:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o6_icb_cmd_sel
                           , o5_icb_cmd_sel
                           , o4_icb_cmd_sel
                           , o3_icb_cmd_sel
                           , o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o6_icb_cmd_valid
                           , o5_icb_cmd_valid
                           , o4_icb_cmd_valid
                           , o3_icb_cmd_valid
                           , o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o6_icb_cmd_read
                           , o5_icb_cmd_read
                           , o4_icb_cmd_read
                           , o3_icb_cmd_read
                           , o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o6_icb_cmd_addr
                           , o5_icb_cmd_addr
                           , o4_icb_cmd_addr
                           , o3_icb_cmd_addr
                           , o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o6_icb_cmd_wdata
                           , o5_icb_cmd_wdata
                           , o4_icb_cmd_wdata
                           , o3_icb_cmd_wdata
                           , o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o6_icb_cmd_wmask
                           , o5_icb_cmd_wmask
                           , o4_icb_cmd_wmask
                           , o3_icb_cmd_wmask
                           , o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o6_icb_cmd_size
                           , o5_icb_cmd_size
                           , o4_icb_cmd_size
                           , o3_icb_cmd_size
                           , o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o6_icb_cmd_lock
                           , o5_icb_cmd_lock
                           , o4_icb_cmd_lock
                           , o3_icb_cmd_lock
                           , o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o6_icb_cmd_excl
                           , o5_icb_cmd_excl
                           , o4_icb_cmd_excl
                           , o3_icb_cmd_excl
                           , o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o6_icb_cmd_xlen
                           , o5_icb_cmd_xlen
                           , o4_icb_cmd_xlen
                           , o3_icb_cmd_xlen
                           , o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o6_icb_cmd_xburst
                           , o5_icb_cmd_xburst
                           , o4_icb_cmd_xburst
                           , o3_icb_cmd_xburst
                           , o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o6_icb_cmd_modes
                           , o5_icb_cmd_modes
                           , o4_icb_cmd_modes
                           , o3_icb_cmd_modes
                           , o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o6_icb_cmd_dmode
                           , o5_icb_cmd_dmode
                           , o4_icb_cmd_dmode
                           , o3_icb_cmd_dmode
                           , o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o6_icb_cmd_attri
                           , o5_icb_cmd_attri
                           , o4_icb_cmd_attri
                           , o3_icb_cmd_attri
                           , o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o6_icb_cmd_beat
                           , o5_icb_cmd_beat
                           , o4_icb_cmd_beat
                           , o3_icb_cmd_beat
                           , o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o6_icb_cmd_usr
                           , o5_icb_cmd_usr
                           , o4_icb_cmd_usr
                           , o3_icb_cmd_usr
                           , o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o6_icb_cmd_ready
                           , o5_icb_cmd_ready
                           , o4_icb_cmd_ready
                           , o3_icb_cmd_ready
                           , o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o6_icb_rsp_valid
                           , o5_icb_rsp_valid
                           , o4_icb_rsp_valid
                           , o3_icb_rsp_valid
                           , o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o6_icb_rsp_err
                           , o5_icb_rsp_err
                           , o4_icb_rsp_err
                           , o3_icb_rsp_err
                           , o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o6_icb_rsp_excl_ok
                           , o5_icb_rsp_excl_ok
                           , o4_icb_rsp_excl_ok
                           , o3_icb_rsp_excl_ok
                           , o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o6_icb_rsp_rdata
                           , o5_icb_rsp_rdata
                           , o4_icb_rsp_rdata
                           , o3_icb_rsp_rdata
                           , o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o6_icb_rsp_usr
                           , o5_icb_rsp_usr
                           , o4_icb_rsp_usr
                           , o3_icb_rsp_usr
                           , o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o6_icb_rsp_ready
                           , o5_icb_rsp_ready
                           , o4_icb_rsp_ready
                           , o3_icb_rsp_ready
                           , o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = (buf_icb_cmd_addr     [31:O2_BASE_REGION_LSB]
                         ==  O2_BASE_ADDR [31:O2_BASE_REGION_LSB] 
                        ) & o2_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
      wire icb_cmd_o3 = (buf_icb_cmd_addr     [31:O3_BASE_REGION_LSB]
                         ==  O3_BASE_ADDR [31:O3_BASE_REGION_LSB] 
                        ) & o3_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                        ; 
      wire icb_cmd_o4 = (buf_icb_cmd_addr     [31:O4_BASE_REGION_LSB]
                         ==  O4_BASE_ADDR [31:O4_BASE_REGION_LSB] 
                        ) & o4_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                        ; 
      wire icb_cmd_o5 = (buf_icb_cmd_addr     [31:O5_BASE_REGION_LSB]
                         ==  O5_BASE_ADDR [31:O5_BASE_REGION_LSB] 
                        ) & o5_icb_enable 
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                        ; 
      wire icb_cmd_o6 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                          & (~icb_cmd_o2)
                          & (~icb_cmd_o3)
                          & (~icb_cmd_o4)
                          & (~icb_cmd_o5)
                        ; 
  wire [7-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o6
                    , icb_cmd_o5
                    , icb_cmd_o4
                    , icb_cmd_o3
                    , icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (7),
  .SPLT_PTR_W (7),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .o_bus_icb_rsp_rdata({(64*7){1'b0}}),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   6:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   6:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   6:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   6:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [ 223:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 447:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  55:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [  20:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   6:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   6:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  55:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [  13:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [  13:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   6:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [  20:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [  13:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [  20:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   6:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   6:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   6:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   6:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [  20:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv0_ro_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (6'b1),
    .i_bus_icb_cmd_wdata({(64*6){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*6)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv1_ro_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (6'b1),
    .i_bus_icb_cmd_wdata({(64*6){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*6)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv2_ro_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (6'b1),
    .i_bus_icb_cmd_wdata({(64*6){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*6)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv3_ro_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (6'b1),
    .i_bus_icb_cmd_wdata({(64*6){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*6)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv4_ro_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (6'b1),
    .i_bus_icb_cmd_wdata({(64*6){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*6)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv5_ro_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (6'b1),
    .i_bus_icb_cmd_wdata({(64*6){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*6)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv6_ro_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (6'b1),
    .i_bus_icb_cmd_wdata({(64*6){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*6)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv0_wo_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (6'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 383:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  47:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv1_wo_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (6'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 383:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  47:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv2_wo_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (6'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 383:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  47:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv3_wo_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (6'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 383:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  47:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv4_wo_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (6'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 383:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  47:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv5_wo_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (6'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 383:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  47:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv6_wo_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire    [   5:   0] arbt_bus_icb_cmd_valid        ;
  wire    [   5:   0] arbt_bus_icb_cmd_ready        ;
  wire    [   5:   0] arbt_bus_icb_cmd_sel          ;
  wire    [   5:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 191:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  47:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  17:   0] arbt_bus_icb_cmd_size         ;
  wire    [   5:   0] arbt_bus_icb_cmd_lock         ;
  wire    [   5:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  47:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  11:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  11:   0] arbt_bus_icb_cmd_modes        ;
  wire    [   5:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  17:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  11:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  17:   0] arbt_bus_icb_cmd_usr          ;
  wire    [   5:   0] arbt_bus_icb_rsp_ready        ;
  wire    [   5:   0] arbt_bus_icb_rsp_valid        ;
  wire    [   5:   0] arbt_bus_icb_rsp_err          ;
  wire    [   5:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 383:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  17:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (6),
  .ARBT_PTR_W (3),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (6'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [   5:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [   5:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 191:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 383:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  47:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  17:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [   5:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [   5:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  47:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  11:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  11:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [   5:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  17:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  11:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  17:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [   5:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [   5:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [   5:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [   5:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 383:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  17:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv0_rw_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
    input              i6_icb_cmd_valid              ,
  output             i6_icb_cmd_ready              ,
  input              i6_icb_cmd_sel                ,
  input              i6_icb_cmd_read               ,
  input  [  31:   0] i6_icb_cmd_addr               ,
  input  [  63:   0] i6_icb_cmd_wdata              ,
  input  [   7:   0] i6_icb_cmd_wmask              ,
  input  [   2:   0] i6_icb_cmd_size               ,
  input              i6_icb_cmd_lock               ,
  input              i6_icb_cmd_excl               ,
  input  [   7:   0] i6_icb_cmd_xlen               ,
  input  [   1:   0] i6_icb_cmd_xburst             ,
  input  [   1:   0] i6_icb_cmd_modes              ,
  input              i6_icb_cmd_dmode              ,
  input  [   2:   0] i6_icb_cmd_attri              ,
  input  [   1:   0] i6_icb_cmd_beat               ,
  input  [   2:   0] i6_icb_cmd_usr                ,
  input              i6_icb_rsp_ready              ,
  output             i6_icb_rsp_valid              ,
  output             i6_icb_rsp_err                ,
  output             i6_icb_rsp_excl_ok            ,
  output [  63:   0] i6_icb_rsp_rdata              ,
  output [   2:   0] i6_icb_rsp_usr                ,
    input              i7_icb_cmd_valid              ,
  output             i7_icb_cmd_ready              ,
  input              i7_icb_cmd_sel                ,
  input              i7_icb_cmd_read               ,
  input  [  31:   0] i7_icb_cmd_addr               ,
  input  [  63:   0] i7_icb_cmd_wdata              ,
  input  [   7:   0] i7_icb_cmd_wmask              ,
  input  [   2:   0] i7_icb_cmd_size               ,
  input              i7_icb_cmd_lock               ,
  input              i7_icb_cmd_excl               ,
  input  [   7:   0] i7_icb_cmd_xlen               ,
  input  [   1:   0] i7_icb_cmd_xburst             ,
  input  [   1:   0] i7_icb_cmd_modes              ,
  input              i7_icb_cmd_dmode              ,
  input  [   2:   0] i7_icb_cmd_attri              ,
  input  [   1:   0] i7_icb_cmd_beat               ,
  input  [   2:   0] i7_icb_cmd_usr                ,
  input              i7_icb_rsp_ready              ,
  output             i7_icb_rsp_valid              ,
  output             i7_icb_rsp_err                ,
  output             i7_icb_rsp_excl_ok            ,
  output [  63:   0] i7_icb_rsp_rdata              ,
  output [   2:   0] i7_icb_rsp_usr                ,
    input              i8_icb_cmd_valid              ,
  output             i8_icb_cmd_ready              ,
  input              i8_icb_cmd_sel                ,
  input              i8_icb_cmd_read               ,
  input  [  31:   0] i8_icb_cmd_addr               ,
  input  [  63:   0] i8_icb_cmd_wdata              ,
  input  [   7:   0] i8_icb_cmd_wmask              ,
  input  [   2:   0] i8_icb_cmd_size               ,
  input              i8_icb_cmd_lock               ,
  input              i8_icb_cmd_excl               ,
  input  [   7:   0] i8_icb_cmd_xlen               ,
  input  [   1:   0] i8_icb_cmd_xburst             ,
  input  [   1:   0] i8_icb_cmd_modes              ,
  input              i8_icb_cmd_dmode              ,
  input  [   2:   0] i8_icb_cmd_attri              ,
  input  [   1:   0] i8_icb_cmd_beat               ,
  input  [   2:   0] i8_icb_cmd_usr                ,
  input              i8_icb_rsp_ready              ,
  output             i8_icb_rsp_valid              ,
  output             i8_icb_rsp_err                ,
  output             i8_icb_rsp_excl_ok            ,
  output [  63:   0] i8_icb_rsp_rdata              ,
  output [   2:   0] i8_icb_rsp_usr                ,
    input              i9_icb_cmd_valid              ,
  output             i9_icb_cmd_ready              ,
  input              i9_icb_cmd_sel                ,
  input              i9_icb_cmd_read               ,
  input  [  31:   0] i9_icb_cmd_addr               ,
  input  [  63:   0] i9_icb_cmd_wdata              ,
  input  [   7:   0] i9_icb_cmd_wmask              ,
  input  [   2:   0] i9_icb_cmd_size               ,
  input              i9_icb_cmd_lock               ,
  input              i9_icb_cmd_excl               ,
  input  [   7:   0] i9_icb_cmd_xlen               ,
  input  [   1:   0] i9_icb_cmd_xburst             ,
  input  [   1:   0] i9_icb_cmd_modes              ,
  input              i9_icb_cmd_dmode              ,
  input  [   2:   0] i9_icb_cmd_attri              ,
  input  [   1:   0] i9_icb_cmd_beat               ,
  input  [   2:   0] i9_icb_cmd_usr                ,
  input              i9_icb_rsp_ready              ,
  output             i9_icb_rsp_valid              ,
  output             i9_icb_rsp_err                ,
  output             i9_icb_rsp_excl_ok            ,
  output [  63:   0] i9_icb_rsp_rdata              ,
  output [   2:   0] i9_icb_rsp_usr                ,
    input              i10_icb_cmd_valid             ,
  output             i10_icb_cmd_ready             ,
  input              i10_icb_cmd_sel               ,
  input              i10_icb_cmd_read              ,
  input  [  31:   0] i10_icb_cmd_addr              ,
  input  [  63:   0] i10_icb_cmd_wdata             ,
  input  [   7:   0] i10_icb_cmd_wmask             ,
  input  [   2:   0] i10_icb_cmd_size              ,
  input              i10_icb_cmd_lock              ,
  input              i10_icb_cmd_excl              ,
  input  [   7:   0] i10_icb_cmd_xlen              ,
  input  [   1:   0] i10_icb_cmd_xburst            ,
  input  [   1:   0] i10_icb_cmd_modes             ,
  input              i10_icb_cmd_dmode             ,
  input  [   2:   0] i10_icb_cmd_attri             ,
  input  [   1:   0] i10_icb_cmd_beat              ,
  input  [   2:   0] i10_icb_cmd_usr               ,
  input              i10_icb_rsp_ready             ,
  output             i10_icb_rsp_valid             ,
  output             i10_icb_rsp_err               ,
  output             i10_icb_rsp_excl_ok           ,
  output [  63:   0] i10_icb_rsp_rdata             ,
  output [   2:   0] i10_icb_rsp_usr               ,
    input              i11_icb_cmd_valid             ,
  output             i11_icb_cmd_ready             ,
  input              i11_icb_cmd_sel               ,
  input              i11_icb_cmd_read              ,
  input  [  31:   0] i11_icb_cmd_addr              ,
  input  [  63:   0] i11_icb_cmd_wdata             ,
  input  [   7:   0] i11_icb_cmd_wmask             ,
  input  [   2:   0] i11_icb_cmd_size              ,
  input              i11_icb_cmd_lock              ,
  input              i11_icb_cmd_excl              ,
  input  [   7:   0] i11_icb_cmd_xlen              ,
  input  [   1:   0] i11_icb_cmd_xburst            ,
  input  [   1:   0] i11_icb_cmd_modes             ,
  input              i11_icb_cmd_dmode             ,
  input  [   2:   0] i11_icb_cmd_attri             ,
  input  [   1:   0] i11_icb_cmd_beat              ,
  input  [   2:   0] i11_icb_cmd_usr               ,
  input              i11_icb_rsp_ready             ,
  output             i11_icb_rsp_valid             ,
  output             i11_icb_rsp_err               ,
  output             i11_icb_rsp_excl_ok           ,
  output [  63:   0] i11_icb_rsp_rdata             ,
  output [   2:   0] i11_icb_rsp_usr               ,
  input  clk,
  input  rst_n
  );
    wire    [  11:   0] arbt_bus_icb_cmd_valid        ;
  wire    [  11:   0] arbt_bus_icb_cmd_ready        ;
  wire    [  11:   0] arbt_bus_icb_cmd_sel          ;
  wire    [  11:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 767:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  95:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  35:   0] arbt_bus_icb_cmd_size         ;
  wire    [  11:   0] arbt_bus_icb_cmd_lock         ;
  wire    [  11:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  95:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  23:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  23:   0] arbt_bus_icb_cmd_modes        ;
  wire    [  11:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  35:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  23:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  35:   0] arbt_bus_icb_cmd_usr          ;
  wire    [  11:   0] arbt_bus_icb_rsp_ready        ;
  wire    [  11:   0] arbt_bus_icb_rsp_valid        ;
  wire    [  11:   0] arbt_bus_icb_rsp_err          ;
  wire    [  11:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 767:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  35:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i11_icb_cmd_valid
                           , i10_icb_cmd_valid
                           , i9_icb_cmd_valid
                           , i8_icb_cmd_valid
                           , i7_icb_cmd_valid
                           , i6_icb_cmd_valid
                           , i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i11_icb_cmd_sel
                           , i10_icb_cmd_sel
                           , i9_icb_cmd_sel
                           , i8_icb_cmd_sel
                           , i7_icb_cmd_sel
                           , i6_icb_cmd_sel
                           , i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i11_icb_cmd_read
                           , i10_icb_cmd_read
                           , i9_icb_cmd_read
                           , i8_icb_cmd_read
                           , i7_icb_cmd_read
                           , i6_icb_cmd_read
                           , i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i11_icb_cmd_addr
                           , i10_icb_cmd_addr
                           , i9_icb_cmd_addr
                           , i8_icb_cmd_addr
                           , i7_icb_cmd_addr
                           , i6_icb_cmd_addr
                           , i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i11_icb_cmd_wdata
                           , i10_icb_cmd_wdata
                           , i9_icb_cmd_wdata
                           , i8_icb_cmd_wdata
                           , i7_icb_cmd_wdata
                           , i6_icb_cmd_wdata
                           , i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i11_icb_cmd_wmask
                           , i10_icb_cmd_wmask
                           , i9_icb_cmd_wmask
                           , i8_icb_cmd_wmask
                           , i7_icb_cmd_wmask
                           , i6_icb_cmd_wmask
                           , i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i11_icb_cmd_size
                           , i10_icb_cmd_size
                           , i9_icb_cmd_size
                           , i8_icb_cmd_size
                           , i7_icb_cmd_size
                           , i6_icb_cmd_size
                           , i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i11_icb_cmd_lock
                           , i10_icb_cmd_lock
                           , i9_icb_cmd_lock
                           , i8_icb_cmd_lock
                           , i7_icb_cmd_lock
                           , i6_icb_cmd_lock
                           , i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i11_icb_cmd_excl
                           , i10_icb_cmd_excl
                           , i9_icb_cmd_excl
                           , i8_icb_cmd_excl
                           , i7_icb_cmd_excl
                           , i6_icb_cmd_excl
                           , i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i11_icb_cmd_xlen
                           , i10_icb_cmd_xlen
                           , i9_icb_cmd_xlen
                           , i8_icb_cmd_xlen
                           , i7_icb_cmd_xlen
                           , i6_icb_cmd_xlen
                           , i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i11_icb_cmd_xburst
                           , i10_icb_cmd_xburst
                           , i9_icb_cmd_xburst
                           , i8_icb_cmd_xburst
                           , i7_icb_cmd_xburst
                           , i6_icb_cmd_xburst
                           , i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i11_icb_cmd_modes
                           , i10_icb_cmd_modes
                           , i9_icb_cmd_modes
                           , i8_icb_cmd_modes
                           , i7_icb_cmd_modes
                           , i6_icb_cmd_modes
                           , i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i11_icb_cmd_dmode
                           , i10_icb_cmd_dmode
                           , i9_icb_cmd_dmode
                           , i8_icb_cmd_dmode
                           , i7_icb_cmd_dmode
                           , i6_icb_cmd_dmode
                           , i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i11_icb_cmd_attri
                           , i10_icb_cmd_attri
                           , i9_icb_cmd_attri
                           , i8_icb_cmd_attri
                           , i7_icb_cmd_attri
                           , i6_icb_cmd_attri
                           , i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i11_icb_cmd_beat
                           , i10_icb_cmd_beat
                           , i9_icb_cmd_beat
                           , i8_icb_cmd_beat
                           , i7_icb_cmd_beat
                           , i6_icb_cmd_beat
                           , i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i11_icb_cmd_usr
                           , i10_icb_cmd_usr
                           , i9_icb_cmd_usr
                           , i8_icb_cmd_usr
                           , i7_icb_cmd_usr
                           , i6_icb_cmd_usr
                           , i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i11_icb_cmd_ready
                           , i10_icb_cmd_ready
                           , i9_icb_cmd_ready
                           , i8_icb_cmd_ready
                           , i7_icb_cmd_ready
                           , i6_icb_cmd_ready
                           , i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i11_icb_rsp_valid
                           , i10_icb_rsp_valid
                           , i9_icb_rsp_valid
                           , i8_icb_rsp_valid
                           , i7_icb_rsp_valid
                           , i6_icb_rsp_valid
                           , i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i11_icb_rsp_err
                           , i10_icb_rsp_err
                           , i9_icb_rsp_err
                           , i8_icb_rsp_err
                           , i7_icb_rsp_err
                           , i6_icb_rsp_err
                           , i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i11_icb_rsp_excl_ok
                           , i10_icb_rsp_excl_ok
                           , i9_icb_rsp_excl_ok
                           , i8_icb_rsp_excl_ok
                           , i7_icb_rsp_excl_ok
                           , i6_icb_rsp_excl_ok
                           , i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i11_icb_rsp_rdata
                           , i10_icb_rsp_rdata
                           , i9_icb_rsp_rdata
                           , i8_icb_rsp_rdata
                           , i7_icb_rsp_rdata
                           , i6_icb_rsp_rdata
                           , i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i11_icb_rsp_usr
                           , i10_icb_rsp_usr
                           , i9_icb_rsp_usr
                           , i8_icb_rsp_usr
                           , i7_icb_rsp_usr
                           , i6_icb_rsp_usr
                           , i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i11_icb_rsp_ready
                           , i10_icb_rsp_ready
                           , i9_icb_rsp_ready
                           , i8_icb_rsp_ready
                           , i7_icb_rsp_ready
                           , i6_icb_rsp_ready
                           , i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (12),
  .ARBT_PTR_W (4),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [  11:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [  11:   0]),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read         [  11:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 383:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 767:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  95:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  35:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [  11:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [  11:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  95:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  23:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  23:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [  11:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  35:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  23:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  35:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [  11:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [  11:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [  11:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [  11:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 767:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  35:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv1_rw_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
    input              i6_icb_cmd_valid              ,
  output             i6_icb_cmd_ready              ,
  input              i6_icb_cmd_sel                ,
  input              i6_icb_cmd_read               ,
  input  [  31:   0] i6_icb_cmd_addr               ,
  input  [  63:   0] i6_icb_cmd_wdata              ,
  input  [   7:   0] i6_icb_cmd_wmask              ,
  input  [   2:   0] i6_icb_cmd_size               ,
  input              i6_icb_cmd_lock               ,
  input              i6_icb_cmd_excl               ,
  input  [   7:   0] i6_icb_cmd_xlen               ,
  input  [   1:   0] i6_icb_cmd_xburst             ,
  input  [   1:   0] i6_icb_cmd_modes              ,
  input              i6_icb_cmd_dmode              ,
  input  [   2:   0] i6_icb_cmd_attri              ,
  input  [   1:   0] i6_icb_cmd_beat               ,
  input  [   2:   0] i6_icb_cmd_usr                ,
  input              i6_icb_rsp_ready              ,
  output             i6_icb_rsp_valid              ,
  output             i6_icb_rsp_err                ,
  output             i6_icb_rsp_excl_ok            ,
  output [  63:   0] i6_icb_rsp_rdata              ,
  output [   2:   0] i6_icb_rsp_usr                ,
    input              i7_icb_cmd_valid              ,
  output             i7_icb_cmd_ready              ,
  input              i7_icb_cmd_sel                ,
  input              i7_icb_cmd_read               ,
  input  [  31:   0] i7_icb_cmd_addr               ,
  input  [  63:   0] i7_icb_cmd_wdata              ,
  input  [   7:   0] i7_icb_cmd_wmask              ,
  input  [   2:   0] i7_icb_cmd_size               ,
  input              i7_icb_cmd_lock               ,
  input              i7_icb_cmd_excl               ,
  input  [   7:   0] i7_icb_cmd_xlen               ,
  input  [   1:   0] i7_icb_cmd_xburst             ,
  input  [   1:   0] i7_icb_cmd_modes              ,
  input              i7_icb_cmd_dmode              ,
  input  [   2:   0] i7_icb_cmd_attri              ,
  input  [   1:   0] i7_icb_cmd_beat               ,
  input  [   2:   0] i7_icb_cmd_usr                ,
  input              i7_icb_rsp_ready              ,
  output             i7_icb_rsp_valid              ,
  output             i7_icb_rsp_err                ,
  output             i7_icb_rsp_excl_ok            ,
  output [  63:   0] i7_icb_rsp_rdata              ,
  output [   2:   0] i7_icb_rsp_usr                ,
    input              i8_icb_cmd_valid              ,
  output             i8_icb_cmd_ready              ,
  input              i8_icb_cmd_sel                ,
  input              i8_icb_cmd_read               ,
  input  [  31:   0] i8_icb_cmd_addr               ,
  input  [  63:   0] i8_icb_cmd_wdata              ,
  input  [   7:   0] i8_icb_cmd_wmask              ,
  input  [   2:   0] i8_icb_cmd_size               ,
  input              i8_icb_cmd_lock               ,
  input              i8_icb_cmd_excl               ,
  input  [   7:   0] i8_icb_cmd_xlen               ,
  input  [   1:   0] i8_icb_cmd_xburst             ,
  input  [   1:   0] i8_icb_cmd_modes              ,
  input              i8_icb_cmd_dmode              ,
  input  [   2:   0] i8_icb_cmd_attri              ,
  input  [   1:   0] i8_icb_cmd_beat               ,
  input  [   2:   0] i8_icb_cmd_usr                ,
  input              i8_icb_rsp_ready              ,
  output             i8_icb_rsp_valid              ,
  output             i8_icb_rsp_err                ,
  output             i8_icb_rsp_excl_ok            ,
  output [  63:   0] i8_icb_rsp_rdata              ,
  output [   2:   0] i8_icb_rsp_usr                ,
    input              i9_icb_cmd_valid              ,
  output             i9_icb_cmd_ready              ,
  input              i9_icb_cmd_sel                ,
  input              i9_icb_cmd_read               ,
  input  [  31:   0] i9_icb_cmd_addr               ,
  input  [  63:   0] i9_icb_cmd_wdata              ,
  input  [   7:   0] i9_icb_cmd_wmask              ,
  input  [   2:   0] i9_icb_cmd_size               ,
  input              i9_icb_cmd_lock               ,
  input              i9_icb_cmd_excl               ,
  input  [   7:   0] i9_icb_cmd_xlen               ,
  input  [   1:   0] i9_icb_cmd_xburst             ,
  input  [   1:   0] i9_icb_cmd_modes              ,
  input              i9_icb_cmd_dmode              ,
  input  [   2:   0] i9_icb_cmd_attri              ,
  input  [   1:   0] i9_icb_cmd_beat               ,
  input  [   2:   0] i9_icb_cmd_usr                ,
  input              i9_icb_rsp_ready              ,
  output             i9_icb_rsp_valid              ,
  output             i9_icb_rsp_err                ,
  output             i9_icb_rsp_excl_ok            ,
  output [  63:   0] i9_icb_rsp_rdata              ,
  output [   2:   0] i9_icb_rsp_usr                ,
    input              i10_icb_cmd_valid             ,
  output             i10_icb_cmd_ready             ,
  input              i10_icb_cmd_sel               ,
  input              i10_icb_cmd_read              ,
  input  [  31:   0] i10_icb_cmd_addr              ,
  input  [  63:   0] i10_icb_cmd_wdata             ,
  input  [   7:   0] i10_icb_cmd_wmask             ,
  input  [   2:   0] i10_icb_cmd_size              ,
  input              i10_icb_cmd_lock              ,
  input              i10_icb_cmd_excl              ,
  input  [   7:   0] i10_icb_cmd_xlen              ,
  input  [   1:   0] i10_icb_cmd_xburst            ,
  input  [   1:   0] i10_icb_cmd_modes             ,
  input              i10_icb_cmd_dmode             ,
  input  [   2:   0] i10_icb_cmd_attri             ,
  input  [   1:   0] i10_icb_cmd_beat              ,
  input  [   2:   0] i10_icb_cmd_usr               ,
  input              i10_icb_rsp_ready             ,
  output             i10_icb_rsp_valid             ,
  output             i10_icb_rsp_err               ,
  output             i10_icb_rsp_excl_ok           ,
  output [  63:   0] i10_icb_rsp_rdata             ,
  output [   2:   0] i10_icb_rsp_usr               ,
    input              i11_icb_cmd_valid             ,
  output             i11_icb_cmd_ready             ,
  input              i11_icb_cmd_sel               ,
  input              i11_icb_cmd_read              ,
  input  [  31:   0] i11_icb_cmd_addr              ,
  input  [  63:   0] i11_icb_cmd_wdata             ,
  input  [   7:   0] i11_icb_cmd_wmask             ,
  input  [   2:   0] i11_icb_cmd_size              ,
  input              i11_icb_cmd_lock              ,
  input              i11_icb_cmd_excl              ,
  input  [   7:   0] i11_icb_cmd_xlen              ,
  input  [   1:   0] i11_icb_cmd_xburst            ,
  input  [   1:   0] i11_icb_cmd_modes             ,
  input              i11_icb_cmd_dmode             ,
  input  [   2:   0] i11_icb_cmd_attri             ,
  input  [   1:   0] i11_icb_cmd_beat              ,
  input  [   2:   0] i11_icb_cmd_usr               ,
  input              i11_icb_rsp_ready             ,
  output             i11_icb_rsp_valid             ,
  output             i11_icb_rsp_err               ,
  output             i11_icb_rsp_excl_ok           ,
  output [  63:   0] i11_icb_rsp_rdata             ,
  output [   2:   0] i11_icb_rsp_usr               ,
  input  clk,
  input  rst_n
  );
    wire    [  11:   0] arbt_bus_icb_cmd_valid        ;
  wire    [  11:   0] arbt_bus_icb_cmd_ready        ;
  wire    [  11:   0] arbt_bus_icb_cmd_sel          ;
  wire    [  11:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 767:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  95:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  35:   0] arbt_bus_icb_cmd_size         ;
  wire    [  11:   0] arbt_bus_icb_cmd_lock         ;
  wire    [  11:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  95:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  23:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  23:   0] arbt_bus_icb_cmd_modes        ;
  wire    [  11:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  35:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  23:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  35:   0] arbt_bus_icb_cmd_usr          ;
  wire    [  11:   0] arbt_bus_icb_rsp_ready        ;
  wire    [  11:   0] arbt_bus_icb_rsp_valid        ;
  wire    [  11:   0] arbt_bus_icb_rsp_err          ;
  wire    [  11:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 767:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  35:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i11_icb_cmd_valid
                           , i10_icb_cmd_valid
                           , i9_icb_cmd_valid
                           , i8_icb_cmd_valid
                           , i7_icb_cmd_valid
                           , i6_icb_cmd_valid
                           , i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i11_icb_cmd_sel
                           , i10_icb_cmd_sel
                           , i9_icb_cmd_sel
                           , i8_icb_cmd_sel
                           , i7_icb_cmd_sel
                           , i6_icb_cmd_sel
                           , i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i11_icb_cmd_read
                           , i10_icb_cmd_read
                           , i9_icb_cmd_read
                           , i8_icb_cmd_read
                           , i7_icb_cmd_read
                           , i6_icb_cmd_read
                           , i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i11_icb_cmd_addr
                           , i10_icb_cmd_addr
                           , i9_icb_cmd_addr
                           , i8_icb_cmd_addr
                           , i7_icb_cmd_addr
                           , i6_icb_cmd_addr
                           , i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i11_icb_cmd_wdata
                           , i10_icb_cmd_wdata
                           , i9_icb_cmd_wdata
                           , i8_icb_cmd_wdata
                           , i7_icb_cmd_wdata
                           , i6_icb_cmd_wdata
                           , i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i11_icb_cmd_wmask
                           , i10_icb_cmd_wmask
                           , i9_icb_cmd_wmask
                           , i8_icb_cmd_wmask
                           , i7_icb_cmd_wmask
                           , i6_icb_cmd_wmask
                           , i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i11_icb_cmd_size
                           , i10_icb_cmd_size
                           , i9_icb_cmd_size
                           , i8_icb_cmd_size
                           , i7_icb_cmd_size
                           , i6_icb_cmd_size
                           , i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i11_icb_cmd_lock
                           , i10_icb_cmd_lock
                           , i9_icb_cmd_lock
                           , i8_icb_cmd_lock
                           , i7_icb_cmd_lock
                           , i6_icb_cmd_lock
                           , i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i11_icb_cmd_excl
                           , i10_icb_cmd_excl
                           , i9_icb_cmd_excl
                           , i8_icb_cmd_excl
                           , i7_icb_cmd_excl
                           , i6_icb_cmd_excl
                           , i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i11_icb_cmd_xlen
                           , i10_icb_cmd_xlen
                           , i9_icb_cmd_xlen
                           , i8_icb_cmd_xlen
                           , i7_icb_cmd_xlen
                           , i6_icb_cmd_xlen
                           , i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i11_icb_cmd_xburst
                           , i10_icb_cmd_xburst
                           , i9_icb_cmd_xburst
                           , i8_icb_cmd_xburst
                           , i7_icb_cmd_xburst
                           , i6_icb_cmd_xburst
                           , i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i11_icb_cmd_modes
                           , i10_icb_cmd_modes
                           , i9_icb_cmd_modes
                           , i8_icb_cmd_modes
                           , i7_icb_cmd_modes
                           , i6_icb_cmd_modes
                           , i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i11_icb_cmd_dmode
                           , i10_icb_cmd_dmode
                           , i9_icb_cmd_dmode
                           , i8_icb_cmd_dmode
                           , i7_icb_cmd_dmode
                           , i6_icb_cmd_dmode
                           , i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i11_icb_cmd_attri
                           , i10_icb_cmd_attri
                           , i9_icb_cmd_attri
                           , i8_icb_cmd_attri
                           , i7_icb_cmd_attri
                           , i6_icb_cmd_attri
                           , i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i11_icb_cmd_beat
                           , i10_icb_cmd_beat
                           , i9_icb_cmd_beat
                           , i8_icb_cmd_beat
                           , i7_icb_cmd_beat
                           , i6_icb_cmd_beat
                           , i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i11_icb_cmd_usr
                           , i10_icb_cmd_usr
                           , i9_icb_cmd_usr
                           , i8_icb_cmd_usr
                           , i7_icb_cmd_usr
                           , i6_icb_cmd_usr
                           , i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i11_icb_cmd_ready
                           , i10_icb_cmd_ready
                           , i9_icb_cmd_ready
                           , i8_icb_cmd_ready
                           , i7_icb_cmd_ready
                           , i6_icb_cmd_ready
                           , i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i11_icb_rsp_valid
                           , i10_icb_rsp_valid
                           , i9_icb_rsp_valid
                           , i8_icb_rsp_valid
                           , i7_icb_rsp_valid
                           , i6_icb_rsp_valid
                           , i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i11_icb_rsp_err
                           , i10_icb_rsp_err
                           , i9_icb_rsp_err
                           , i8_icb_rsp_err
                           , i7_icb_rsp_err
                           , i6_icb_rsp_err
                           , i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i11_icb_rsp_excl_ok
                           , i10_icb_rsp_excl_ok
                           , i9_icb_rsp_excl_ok
                           , i8_icb_rsp_excl_ok
                           , i7_icb_rsp_excl_ok
                           , i6_icb_rsp_excl_ok
                           , i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i11_icb_rsp_rdata
                           , i10_icb_rsp_rdata
                           , i9_icb_rsp_rdata
                           , i8_icb_rsp_rdata
                           , i7_icb_rsp_rdata
                           , i6_icb_rsp_rdata
                           , i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i11_icb_rsp_usr
                           , i10_icb_rsp_usr
                           , i9_icb_rsp_usr
                           , i8_icb_rsp_usr
                           , i7_icb_rsp_usr
                           , i6_icb_rsp_usr
                           , i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i11_icb_rsp_ready
                           , i10_icb_rsp_ready
                           , i9_icb_rsp_ready
                           , i8_icb_rsp_ready
                           , i7_icb_rsp_ready
                           , i6_icb_rsp_ready
                           , i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (12),
  .ARBT_PTR_W (4),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [  11:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [  11:   0]),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read         [  11:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 383:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 767:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  95:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  35:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [  11:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [  11:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  95:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  23:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  23:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [  11:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  35:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  23:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  35:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [  11:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [  11:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [  11:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [  11:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 767:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  35:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv2_rw_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
    input              i6_icb_cmd_valid              ,
  output             i6_icb_cmd_ready              ,
  input              i6_icb_cmd_sel                ,
  input              i6_icb_cmd_read               ,
  input  [  31:   0] i6_icb_cmd_addr               ,
  input  [  63:   0] i6_icb_cmd_wdata              ,
  input  [   7:   0] i6_icb_cmd_wmask              ,
  input  [   2:   0] i6_icb_cmd_size               ,
  input              i6_icb_cmd_lock               ,
  input              i6_icb_cmd_excl               ,
  input  [   7:   0] i6_icb_cmd_xlen               ,
  input  [   1:   0] i6_icb_cmd_xburst             ,
  input  [   1:   0] i6_icb_cmd_modes              ,
  input              i6_icb_cmd_dmode              ,
  input  [   2:   0] i6_icb_cmd_attri              ,
  input  [   1:   0] i6_icb_cmd_beat               ,
  input  [   2:   0] i6_icb_cmd_usr                ,
  input              i6_icb_rsp_ready              ,
  output             i6_icb_rsp_valid              ,
  output             i6_icb_rsp_err                ,
  output             i6_icb_rsp_excl_ok            ,
  output [  63:   0] i6_icb_rsp_rdata              ,
  output [   2:   0] i6_icb_rsp_usr                ,
    input              i7_icb_cmd_valid              ,
  output             i7_icb_cmd_ready              ,
  input              i7_icb_cmd_sel                ,
  input              i7_icb_cmd_read               ,
  input  [  31:   0] i7_icb_cmd_addr               ,
  input  [  63:   0] i7_icb_cmd_wdata              ,
  input  [   7:   0] i7_icb_cmd_wmask              ,
  input  [   2:   0] i7_icb_cmd_size               ,
  input              i7_icb_cmd_lock               ,
  input              i7_icb_cmd_excl               ,
  input  [   7:   0] i7_icb_cmd_xlen               ,
  input  [   1:   0] i7_icb_cmd_xburst             ,
  input  [   1:   0] i7_icb_cmd_modes              ,
  input              i7_icb_cmd_dmode              ,
  input  [   2:   0] i7_icb_cmd_attri              ,
  input  [   1:   0] i7_icb_cmd_beat               ,
  input  [   2:   0] i7_icb_cmd_usr                ,
  input              i7_icb_rsp_ready              ,
  output             i7_icb_rsp_valid              ,
  output             i7_icb_rsp_err                ,
  output             i7_icb_rsp_excl_ok            ,
  output [  63:   0] i7_icb_rsp_rdata              ,
  output [   2:   0] i7_icb_rsp_usr                ,
    input              i8_icb_cmd_valid              ,
  output             i8_icb_cmd_ready              ,
  input              i8_icb_cmd_sel                ,
  input              i8_icb_cmd_read               ,
  input  [  31:   0] i8_icb_cmd_addr               ,
  input  [  63:   0] i8_icb_cmd_wdata              ,
  input  [   7:   0] i8_icb_cmd_wmask              ,
  input  [   2:   0] i8_icb_cmd_size               ,
  input              i8_icb_cmd_lock               ,
  input              i8_icb_cmd_excl               ,
  input  [   7:   0] i8_icb_cmd_xlen               ,
  input  [   1:   0] i8_icb_cmd_xburst             ,
  input  [   1:   0] i8_icb_cmd_modes              ,
  input              i8_icb_cmd_dmode              ,
  input  [   2:   0] i8_icb_cmd_attri              ,
  input  [   1:   0] i8_icb_cmd_beat               ,
  input  [   2:   0] i8_icb_cmd_usr                ,
  input              i8_icb_rsp_ready              ,
  output             i8_icb_rsp_valid              ,
  output             i8_icb_rsp_err                ,
  output             i8_icb_rsp_excl_ok            ,
  output [  63:   0] i8_icb_rsp_rdata              ,
  output [   2:   0] i8_icb_rsp_usr                ,
    input              i9_icb_cmd_valid              ,
  output             i9_icb_cmd_ready              ,
  input              i9_icb_cmd_sel                ,
  input              i9_icb_cmd_read               ,
  input  [  31:   0] i9_icb_cmd_addr               ,
  input  [  63:   0] i9_icb_cmd_wdata              ,
  input  [   7:   0] i9_icb_cmd_wmask              ,
  input  [   2:   0] i9_icb_cmd_size               ,
  input              i9_icb_cmd_lock               ,
  input              i9_icb_cmd_excl               ,
  input  [   7:   0] i9_icb_cmd_xlen               ,
  input  [   1:   0] i9_icb_cmd_xburst             ,
  input  [   1:   0] i9_icb_cmd_modes              ,
  input              i9_icb_cmd_dmode              ,
  input  [   2:   0] i9_icb_cmd_attri              ,
  input  [   1:   0] i9_icb_cmd_beat               ,
  input  [   2:   0] i9_icb_cmd_usr                ,
  input              i9_icb_rsp_ready              ,
  output             i9_icb_rsp_valid              ,
  output             i9_icb_rsp_err                ,
  output             i9_icb_rsp_excl_ok            ,
  output [  63:   0] i9_icb_rsp_rdata              ,
  output [   2:   0] i9_icb_rsp_usr                ,
    input              i10_icb_cmd_valid             ,
  output             i10_icb_cmd_ready             ,
  input              i10_icb_cmd_sel               ,
  input              i10_icb_cmd_read              ,
  input  [  31:   0] i10_icb_cmd_addr              ,
  input  [  63:   0] i10_icb_cmd_wdata             ,
  input  [   7:   0] i10_icb_cmd_wmask             ,
  input  [   2:   0] i10_icb_cmd_size              ,
  input              i10_icb_cmd_lock              ,
  input              i10_icb_cmd_excl              ,
  input  [   7:   0] i10_icb_cmd_xlen              ,
  input  [   1:   0] i10_icb_cmd_xburst            ,
  input  [   1:   0] i10_icb_cmd_modes             ,
  input              i10_icb_cmd_dmode             ,
  input  [   2:   0] i10_icb_cmd_attri             ,
  input  [   1:   0] i10_icb_cmd_beat              ,
  input  [   2:   0] i10_icb_cmd_usr               ,
  input              i10_icb_rsp_ready             ,
  output             i10_icb_rsp_valid             ,
  output             i10_icb_rsp_err               ,
  output             i10_icb_rsp_excl_ok           ,
  output [  63:   0] i10_icb_rsp_rdata             ,
  output [   2:   0] i10_icb_rsp_usr               ,
    input              i11_icb_cmd_valid             ,
  output             i11_icb_cmd_ready             ,
  input              i11_icb_cmd_sel               ,
  input              i11_icb_cmd_read              ,
  input  [  31:   0] i11_icb_cmd_addr              ,
  input  [  63:   0] i11_icb_cmd_wdata             ,
  input  [   7:   0] i11_icb_cmd_wmask             ,
  input  [   2:   0] i11_icb_cmd_size              ,
  input              i11_icb_cmd_lock              ,
  input              i11_icb_cmd_excl              ,
  input  [   7:   0] i11_icb_cmd_xlen              ,
  input  [   1:   0] i11_icb_cmd_xburst            ,
  input  [   1:   0] i11_icb_cmd_modes             ,
  input              i11_icb_cmd_dmode             ,
  input  [   2:   0] i11_icb_cmd_attri             ,
  input  [   1:   0] i11_icb_cmd_beat              ,
  input  [   2:   0] i11_icb_cmd_usr               ,
  input              i11_icb_rsp_ready             ,
  output             i11_icb_rsp_valid             ,
  output             i11_icb_rsp_err               ,
  output             i11_icb_rsp_excl_ok           ,
  output [  63:   0] i11_icb_rsp_rdata             ,
  output [   2:   0] i11_icb_rsp_usr               ,
  input  clk,
  input  rst_n
  );
    wire    [  11:   0] arbt_bus_icb_cmd_valid        ;
  wire    [  11:   0] arbt_bus_icb_cmd_ready        ;
  wire    [  11:   0] arbt_bus_icb_cmd_sel          ;
  wire    [  11:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 767:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  95:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  35:   0] arbt_bus_icb_cmd_size         ;
  wire    [  11:   0] arbt_bus_icb_cmd_lock         ;
  wire    [  11:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  95:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  23:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  23:   0] arbt_bus_icb_cmd_modes        ;
  wire    [  11:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  35:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  23:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  35:   0] arbt_bus_icb_cmd_usr          ;
  wire    [  11:   0] arbt_bus_icb_rsp_ready        ;
  wire    [  11:   0] arbt_bus_icb_rsp_valid        ;
  wire    [  11:   0] arbt_bus_icb_rsp_err          ;
  wire    [  11:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 767:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  35:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i11_icb_cmd_valid
                           , i10_icb_cmd_valid
                           , i9_icb_cmd_valid
                           , i8_icb_cmd_valid
                           , i7_icb_cmd_valid
                           , i6_icb_cmd_valid
                           , i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i11_icb_cmd_sel
                           , i10_icb_cmd_sel
                           , i9_icb_cmd_sel
                           , i8_icb_cmd_sel
                           , i7_icb_cmd_sel
                           , i6_icb_cmd_sel
                           , i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i11_icb_cmd_read
                           , i10_icb_cmd_read
                           , i9_icb_cmd_read
                           , i8_icb_cmd_read
                           , i7_icb_cmd_read
                           , i6_icb_cmd_read
                           , i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i11_icb_cmd_addr
                           , i10_icb_cmd_addr
                           , i9_icb_cmd_addr
                           , i8_icb_cmd_addr
                           , i7_icb_cmd_addr
                           , i6_icb_cmd_addr
                           , i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i11_icb_cmd_wdata
                           , i10_icb_cmd_wdata
                           , i9_icb_cmd_wdata
                           , i8_icb_cmd_wdata
                           , i7_icb_cmd_wdata
                           , i6_icb_cmd_wdata
                           , i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i11_icb_cmd_wmask
                           , i10_icb_cmd_wmask
                           , i9_icb_cmd_wmask
                           , i8_icb_cmd_wmask
                           , i7_icb_cmd_wmask
                           , i6_icb_cmd_wmask
                           , i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i11_icb_cmd_size
                           , i10_icb_cmd_size
                           , i9_icb_cmd_size
                           , i8_icb_cmd_size
                           , i7_icb_cmd_size
                           , i6_icb_cmd_size
                           , i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i11_icb_cmd_lock
                           , i10_icb_cmd_lock
                           , i9_icb_cmd_lock
                           , i8_icb_cmd_lock
                           , i7_icb_cmd_lock
                           , i6_icb_cmd_lock
                           , i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i11_icb_cmd_excl
                           , i10_icb_cmd_excl
                           , i9_icb_cmd_excl
                           , i8_icb_cmd_excl
                           , i7_icb_cmd_excl
                           , i6_icb_cmd_excl
                           , i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i11_icb_cmd_xlen
                           , i10_icb_cmd_xlen
                           , i9_icb_cmd_xlen
                           , i8_icb_cmd_xlen
                           , i7_icb_cmd_xlen
                           , i6_icb_cmd_xlen
                           , i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i11_icb_cmd_xburst
                           , i10_icb_cmd_xburst
                           , i9_icb_cmd_xburst
                           , i8_icb_cmd_xburst
                           , i7_icb_cmd_xburst
                           , i6_icb_cmd_xburst
                           , i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i11_icb_cmd_modes
                           , i10_icb_cmd_modes
                           , i9_icb_cmd_modes
                           , i8_icb_cmd_modes
                           , i7_icb_cmd_modes
                           , i6_icb_cmd_modes
                           , i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i11_icb_cmd_dmode
                           , i10_icb_cmd_dmode
                           , i9_icb_cmd_dmode
                           , i8_icb_cmd_dmode
                           , i7_icb_cmd_dmode
                           , i6_icb_cmd_dmode
                           , i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i11_icb_cmd_attri
                           , i10_icb_cmd_attri
                           , i9_icb_cmd_attri
                           , i8_icb_cmd_attri
                           , i7_icb_cmd_attri
                           , i6_icb_cmd_attri
                           , i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i11_icb_cmd_beat
                           , i10_icb_cmd_beat
                           , i9_icb_cmd_beat
                           , i8_icb_cmd_beat
                           , i7_icb_cmd_beat
                           , i6_icb_cmd_beat
                           , i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i11_icb_cmd_usr
                           , i10_icb_cmd_usr
                           , i9_icb_cmd_usr
                           , i8_icb_cmd_usr
                           , i7_icb_cmd_usr
                           , i6_icb_cmd_usr
                           , i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i11_icb_cmd_ready
                           , i10_icb_cmd_ready
                           , i9_icb_cmd_ready
                           , i8_icb_cmd_ready
                           , i7_icb_cmd_ready
                           , i6_icb_cmd_ready
                           , i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i11_icb_rsp_valid
                           , i10_icb_rsp_valid
                           , i9_icb_rsp_valid
                           , i8_icb_rsp_valid
                           , i7_icb_rsp_valid
                           , i6_icb_rsp_valid
                           , i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i11_icb_rsp_err
                           , i10_icb_rsp_err
                           , i9_icb_rsp_err
                           , i8_icb_rsp_err
                           , i7_icb_rsp_err
                           , i6_icb_rsp_err
                           , i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i11_icb_rsp_excl_ok
                           , i10_icb_rsp_excl_ok
                           , i9_icb_rsp_excl_ok
                           , i8_icb_rsp_excl_ok
                           , i7_icb_rsp_excl_ok
                           , i6_icb_rsp_excl_ok
                           , i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i11_icb_rsp_rdata
                           , i10_icb_rsp_rdata
                           , i9_icb_rsp_rdata
                           , i8_icb_rsp_rdata
                           , i7_icb_rsp_rdata
                           , i6_icb_rsp_rdata
                           , i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i11_icb_rsp_usr
                           , i10_icb_rsp_usr
                           , i9_icb_rsp_usr
                           , i8_icb_rsp_usr
                           , i7_icb_rsp_usr
                           , i6_icb_rsp_usr
                           , i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i11_icb_rsp_ready
                           , i10_icb_rsp_ready
                           , i9_icb_rsp_ready
                           , i8_icb_rsp_ready
                           , i7_icb_rsp_ready
                           , i6_icb_rsp_ready
                           , i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (12),
  .ARBT_PTR_W (4),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [  11:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [  11:   0]),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read         [  11:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 383:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 767:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  95:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  35:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [  11:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [  11:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  95:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  23:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  23:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [  11:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  35:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  23:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  35:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [  11:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [  11:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [  11:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [  11:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 767:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  35:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv3_rw_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
    input              i6_icb_cmd_valid              ,
  output             i6_icb_cmd_ready              ,
  input              i6_icb_cmd_sel                ,
  input              i6_icb_cmd_read               ,
  input  [  31:   0] i6_icb_cmd_addr               ,
  input  [  63:   0] i6_icb_cmd_wdata              ,
  input  [   7:   0] i6_icb_cmd_wmask              ,
  input  [   2:   0] i6_icb_cmd_size               ,
  input              i6_icb_cmd_lock               ,
  input              i6_icb_cmd_excl               ,
  input  [   7:   0] i6_icb_cmd_xlen               ,
  input  [   1:   0] i6_icb_cmd_xburst             ,
  input  [   1:   0] i6_icb_cmd_modes              ,
  input              i6_icb_cmd_dmode              ,
  input  [   2:   0] i6_icb_cmd_attri              ,
  input  [   1:   0] i6_icb_cmd_beat               ,
  input  [   2:   0] i6_icb_cmd_usr                ,
  input              i6_icb_rsp_ready              ,
  output             i6_icb_rsp_valid              ,
  output             i6_icb_rsp_err                ,
  output             i6_icb_rsp_excl_ok            ,
  output [  63:   0] i6_icb_rsp_rdata              ,
  output [   2:   0] i6_icb_rsp_usr                ,
    input              i7_icb_cmd_valid              ,
  output             i7_icb_cmd_ready              ,
  input              i7_icb_cmd_sel                ,
  input              i7_icb_cmd_read               ,
  input  [  31:   0] i7_icb_cmd_addr               ,
  input  [  63:   0] i7_icb_cmd_wdata              ,
  input  [   7:   0] i7_icb_cmd_wmask              ,
  input  [   2:   0] i7_icb_cmd_size               ,
  input              i7_icb_cmd_lock               ,
  input              i7_icb_cmd_excl               ,
  input  [   7:   0] i7_icb_cmd_xlen               ,
  input  [   1:   0] i7_icb_cmd_xburst             ,
  input  [   1:   0] i7_icb_cmd_modes              ,
  input              i7_icb_cmd_dmode              ,
  input  [   2:   0] i7_icb_cmd_attri              ,
  input  [   1:   0] i7_icb_cmd_beat               ,
  input  [   2:   0] i7_icb_cmd_usr                ,
  input              i7_icb_rsp_ready              ,
  output             i7_icb_rsp_valid              ,
  output             i7_icb_rsp_err                ,
  output             i7_icb_rsp_excl_ok            ,
  output [  63:   0] i7_icb_rsp_rdata              ,
  output [   2:   0] i7_icb_rsp_usr                ,
    input              i8_icb_cmd_valid              ,
  output             i8_icb_cmd_ready              ,
  input              i8_icb_cmd_sel                ,
  input              i8_icb_cmd_read               ,
  input  [  31:   0] i8_icb_cmd_addr               ,
  input  [  63:   0] i8_icb_cmd_wdata              ,
  input  [   7:   0] i8_icb_cmd_wmask              ,
  input  [   2:   0] i8_icb_cmd_size               ,
  input              i8_icb_cmd_lock               ,
  input              i8_icb_cmd_excl               ,
  input  [   7:   0] i8_icb_cmd_xlen               ,
  input  [   1:   0] i8_icb_cmd_xburst             ,
  input  [   1:   0] i8_icb_cmd_modes              ,
  input              i8_icb_cmd_dmode              ,
  input  [   2:   0] i8_icb_cmd_attri              ,
  input  [   1:   0] i8_icb_cmd_beat               ,
  input  [   2:   0] i8_icb_cmd_usr                ,
  input              i8_icb_rsp_ready              ,
  output             i8_icb_rsp_valid              ,
  output             i8_icb_rsp_err                ,
  output             i8_icb_rsp_excl_ok            ,
  output [  63:   0] i8_icb_rsp_rdata              ,
  output [   2:   0] i8_icb_rsp_usr                ,
    input              i9_icb_cmd_valid              ,
  output             i9_icb_cmd_ready              ,
  input              i9_icb_cmd_sel                ,
  input              i9_icb_cmd_read               ,
  input  [  31:   0] i9_icb_cmd_addr               ,
  input  [  63:   0] i9_icb_cmd_wdata              ,
  input  [   7:   0] i9_icb_cmd_wmask              ,
  input  [   2:   0] i9_icb_cmd_size               ,
  input              i9_icb_cmd_lock               ,
  input              i9_icb_cmd_excl               ,
  input  [   7:   0] i9_icb_cmd_xlen               ,
  input  [   1:   0] i9_icb_cmd_xburst             ,
  input  [   1:   0] i9_icb_cmd_modes              ,
  input              i9_icb_cmd_dmode              ,
  input  [   2:   0] i9_icb_cmd_attri              ,
  input  [   1:   0] i9_icb_cmd_beat               ,
  input  [   2:   0] i9_icb_cmd_usr                ,
  input              i9_icb_rsp_ready              ,
  output             i9_icb_rsp_valid              ,
  output             i9_icb_rsp_err                ,
  output             i9_icb_rsp_excl_ok            ,
  output [  63:   0] i9_icb_rsp_rdata              ,
  output [   2:   0] i9_icb_rsp_usr                ,
    input              i10_icb_cmd_valid             ,
  output             i10_icb_cmd_ready             ,
  input              i10_icb_cmd_sel               ,
  input              i10_icb_cmd_read              ,
  input  [  31:   0] i10_icb_cmd_addr              ,
  input  [  63:   0] i10_icb_cmd_wdata             ,
  input  [   7:   0] i10_icb_cmd_wmask             ,
  input  [   2:   0] i10_icb_cmd_size              ,
  input              i10_icb_cmd_lock              ,
  input              i10_icb_cmd_excl              ,
  input  [   7:   0] i10_icb_cmd_xlen              ,
  input  [   1:   0] i10_icb_cmd_xburst            ,
  input  [   1:   0] i10_icb_cmd_modes             ,
  input              i10_icb_cmd_dmode             ,
  input  [   2:   0] i10_icb_cmd_attri             ,
  input  [   1:   0] i10_icb_cmd_beat              ,
  input  [   2:   0] i10_icb_cmd_usr               ,
  input              i10_icb_rsp_ready             ,
  output             i10_icb_rsp_valid             ,
  output             i10_icb_rsp_err               ,
  output             i10_icb_rsp_excl_ok           ,
  output [  63:   0] i10_icb_rsp_rdata             ,
  output [   2:   0] i10_icb_rsp_usr               ,
    input              i11_icb_cmd_valid             ,
  output             i11_icb_cmd_ready             ,
  input              i11_icb_cmd_sel               ,
  input              i11_icb_cmd_read              ,
  input  [  31:   0] i11_icb_cmd_addr              ,
  input  [  63:   0] i11_icb_cmd_wdata             ,
  input  [   7:   0] i11_icb_cmd_wmask             ,
  input  [   2:   0] i11_icb_cmd_size              ,
  input              i11_icb_cmd_lock              ,
  input              i11_icb_cmd_excl              ,
  input  [   7:   0] i11_icb_cmd_xlen              ,
  input  [   1:   0] i11_icb_cmd_xburst            ,
  input  [   1:   0] i11_icb_cmd_modes             ,
  input              i11_icb_cmd_dmode             ,
  input  [   2:   0] i11_icb_cmd_attri             ,
  input  [   1:   0] i11_icb_cmd_beat              ,
  input  [   2:   0] i11_icb_cmd_usr               ,
  input              i11_icb_rsp_ready             ,
  output             i11_icb_rsp_valid             ,
  output             i11_icb_rsp_err               ,
  output             i11_icb_rsp_excl_ok           ,
  output [  63:   0] i11_icb_rsp_rdata             ,
  output [   2:   0] i11_icb_rsp_usr               ,
  input  clk,
  input  rst_n
  );
    wire    [  11:   0] arbt_bus_icb_cmd_valid        ;
  wire    [  11:   0] arbt_bus_icb_cmd_ready        ;
  wire    [  11:   0] arbt_bus_icb_cmd_sel          ;
  wire    [  11:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 767:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  95:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  35:   0] arbt_bus_icb_cmd_size         ;
  wire    [  11:   0] arbt_bus_icb_cmd_lock         ;
  wire    [  11:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  95:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  23:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  23:   0] arbt_bus_icb_cmd_modes        ;
  wire    [  11:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  35:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  23:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  35:   0] arbt_bus_icb_cmd_usr          ;
  wire    [  11:   0] arbt_bus_icb_rsp_ready        ;
  wire    [  11:   0] arbt_bus_icb_rsp_valid        ;
  wire    [  11:   0] arbt_bus_icb_rsp_err          ;
  wire    [  11:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 767:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  35:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i11_icb_cmd_valid
                           , i10_icb_cmd_valid
                           , i9_icb_cmd_valid
                           , i8_icb_cmd_valid
                           , i7_icb_cmd_valid
                           , i6_icb_cmd_valid
                           , i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i11_icb_cmd_sel
                           , i10_icb_cmd_sel
                           , i9_icb_cmd_sel
                           , i8_icb_cmd_sel
                           , i7_icb_cmd_sel
                           , i6_icb_cmd_sel
                           , i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i11_icb_cmd_read
                           , i10_icb_cmd_read
                           , i9_icb_cmd_read
                           , i8_icb_cmd_read
                           , i7_icb_cmd_read
                           , i6_icb_cmd_read
                           , i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i11_icb_cmd_addr
                           , i10_icb_cmd_addr
                           , i9_icb_cmd_addr
                           , i8_icb_cmd_addr
                           , i7_icb_cmd_addr
                           , i6_icb_cmd_addr
                           , i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i11_icb_cmd_wdata
                           , i10_icb_cmd_wdata
                           , i9_icb_cmd_wdata
                           , i8_icb_cmd_wdata
                           , i7_icb_cmd_wdata
                           , i6_icb_cmd_wdata
                           , i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i11_icb_cmd_wmask
                           , i10_icb_cmd_wmask
                           , i9_icb_cmd_wmask
                           , i8_icb_cmd_wmask
                           , i7_icb_cmd_wmask
                           , i6_icb_cmd_wmask
                           , i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i11_icb_cmd_size
                           , i10_icb_cmd_size
                           , i9_icb_cmd_size
                           , i8_icb_cmd_size
                           , i7_icb_cmd_size
                           , i6_icb_cmd_size
                           , i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i11_icb_cmd_lock
                           , i10_icb_cmd_lock
                           , i9_icb_cmd_lock
                           , i8_icb_cmd_lock
                           , i7_icb_cmd_lock
                           , i6_icb_cmd_lock
                           , i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i11_icb_cmd_excl
                           , i10_icb_cmd_excl
                           , i9_icb_cmd_excl
                           , i8_icb_cmd_excl
                           , i7_icb_cmd_excl
                           , i6_icb_cmd_excl
                           , i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i11_icb_cmd_xlen
                           , i10_icb_cmd_xlen
                           , i9_icb_cmd_xlen
                           , i8_icb_cmd_xlen
                           , i7_icb_cmd_xlen
                           , i6_icb_cmd_xlen
                           , i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i11_icb_cmd_xburst
                           , i10_icb_cmd_xburst
                           , i9_icb_cmd_xburst
                           , i8_icb_cmd_xburst
                           , i7_icb_cmd_xburst
                           , i6_icb_cmd_xburst
                           , i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i11_icb_cmd_modes
                           , i10_icb_cmd_modes
                           , i9_icb_cmd_modes
                           , i8_icb_cmd_modes
                           , i7_icb_cmd_modes
                           , i6_icb_cmd_modes
                           , i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i11_icb_cmd_dmode
                           , i10_icb_cmd_dmode
                           , i9_icb_cmd_dmode
                           , i8_icb_cmd_dmode
                           , i7_icb_cmd_dmode
                           , i6_icb_cmd_dmode
                           , i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i11_icb_cmd_attri
                           , i10_icb_cmd_attri
                           , i9_icb_cmd_attri
                           , i8_icb_cmd_attri
                           , i7_icb_cmd_attri
                           , i6_icb_cmd_attri
                           , i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i11_icb_cmd_beat
                           , i10_icb_cmd_beat
                           , i9_icb_cmd_beat
                           , i8_icb_cmd_beat
                           , i7_icb_cmd_beat
                           , i6_icb_cmd_beat
                           , i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i11_icb_cmd_usr
                           , i10_icb_cmd_usr
                           , i9_icb_cmd_usr
                           , i8_icb_cmd_usr
                           , i7_icb_cmd_usr
                           , i6_icb_cmd_usr
                           , i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i11_icb_cmd_ready
                           , i10_icb_cmd_ready
                           , i9_icb_cmd_ready
                           , i8_icb_cmd_ready
                           , i7_icb_cmd_ready
                           , i6_icb_cmd_ready
                           , i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i11_icb_rsp_valid
                           , i10_icb_rsp_valid
                           , i9_icb_rsp_valid
                           , i8_icb_rsp_valid
                           , i7_icb_rsp_valid
                           , i6_icb_rsp_valid
                           , i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i11_icb_rsp_err
                           , i10_icb_rsp_err
                           , i9_icb_rsp_err
                           , i8_icb_rsp_err
                           , i7_icb_rsp_err
                           , i6_icb_rsp_err
                           , i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i11_icb_rsp_excl_ok
                           , i10_icb_rsp_excl_ok
                           , i9_icb_rsp_excl_ok
                           , i8_icb_rsp_excl_ok
                           , i7_icb_rsp_excl_ok
                           , i6_icb_rsp_excl_ok
                           , i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i11_icb_rsp_rdata
                           , i10_icb_rsp_rdata
                           , i9_icb_rsp_rdata
                           , i8_icb_rsp_rdata
                           , i7_icb_rsp_rdata
                           , i6_icb_rsp_rdata
                           , i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i11_icb_rsp_usr
                           , i10_icb_rsp_usr
                           , i9_icb_rsp_usr
                           , i8_icb_rsp_usr
                           , i7_icb_rsp_usr
                           , i6_icb_rsp_usr
                           , i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i11_icb_rsp_ready
                           , i10_icb_rsp_ready
                           , i9_icb_rsp_ready
                           , i8_icb_rsp_ready
                           , i7_icb_rsp_ready
                           , i6_icb_rsp_ready
                           , i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (12),
  .ARBT_PTR_W (4),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [  11:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [  11:   0]),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read         [  11:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 383:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 767:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  95:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  35:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [  11:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [  11:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  95:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  23:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  23:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [  11:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  35:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  23:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  35:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [  11:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [  11:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [  11:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [  11:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 767:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  35:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv4_rw_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
    input              i6_icb_cmd_valid              ,
  output             i6_icb_cmd_ready              ,
  input              i6_icb_cmd_sel                ,
  input              i6_icb_cmd_read               ,
  input  [  31:   0] i6_icb_cmd_addr               ,
  input  [  63:   0] i6_icb_cmd_wdata              ,
  input  [   7:   0] i6_icb_cmd_wmask              ,
  input  [   2:   0] i6_icb_cmd_size               ,
  input              i6_icb_cmd_lock               ,
  input              i6_icb_cmd_excl               ,
  input  [   7:   0] i6_icb_cmd_xlen               ,
  input  [   1:   0] i6_icb_cmd_xburst             ,
  input  [   1:   0] i6_icb_cmd_modes              ,
  input              i6_icb_cmd_dmode              ,
  input  [   2:   0] i6_icb_cmd_attri              ,
  input  [   1:   0] i6_icb_cmd_beat               ,
  input  [   2:   0] i6_icb_cmd_usr                ,
  input              i6_icb_rsp_ready              ,
  output             i6_icb_rsp_valid              ,
  output             i6_icb_rsp_err                ,
  output             i6_icb_rsp_excl_ok            ,
  output [  63:   0] i6_icb_rsp_rdata              ,
  output [   2:   0] i6_icb_rsp_usr                ,
    input              i7_icb_cmd_valid              ,
  output             i7_icb_cmd_ready              ,
  input              i7_icb_cmd_sel                ,
  input              i7_icb_cmd_read               ,
  input  [  31:   0] i7_icb_cmd_addr               ,
  input  [  63:   0] i7_icb_cmd_wdata              ,
  input  [   7:   0] i7_icb_cmd_wmask              ,
  input  [   2:   0] i7_icb_cmd_size               ,
  input              i7_icb_cmd_lock               ,
  input              i7_icb_cmd_excl               ,
  input  [   7:   0] i7_icb_cmd_xlen               ,
  input  [   1:   0] i7_icb_cmd_xburst             ,
  input  [   1:   0] i7_icb_cmd_modes              ,
  input              i7_icb_cmd_dmode              ,
  input  [   2:   0] i7_icb_cmd_attri              ,
  input  [   1:   0] i7_icb_cmd_beat               ,
  input  [   2:   0] i7_icb_cmd_usr                ,
  input              i7_icb_rsp_ready              ,
  output             i7_icb_rsp_valid              ,
  output             i7_icb_rsp_err                ,
  output             i7_icb_rsp_excl_ok            ,
  output [  63:   0] i7_icb_rsp_rdata              ,
  output [   2:   0] i7_icb_rsp_usr                ,
    input              i8_icb_cmd_valid              ,
  output             i8_icb_cmd_ready              ,
  input              i8_icb_cmd_sel                ,
  input              i8_icb_cmd_read               ,
  input  [  31:   0] i8_icb_cmd_addr               ,
  input  [  63:   0] i8_icb_cmd_wdata              ,
  input  [   7:   0] i8_icb_cmd_wmask              ,
  input  [   2:   0] i8_icb_cmd_size               ,
  input              i8_icb_cmd_lock               ,
  input              i8_icb_cmd_excl               ,
  input  [   7:   0] i8_icb_cmd_xlen               ,
  input  [   1:   0] i8_icb_cmd_xburst             ,
  input  [   1:   0] i8_icb_cmd_modes              ,
  input              i8_icb_cmd_dmode              ,
  input  [   2:   0] i8_icb_cmd_attri              ,
  input  [   1:   0] i8_icb_cmd_beat               ,
  input  [   2:   0] i8_icb_cmd_usr                ,
  input              i8_icb_rsp_ready              ,
  output             i8_icb_rsp_valid              ,
  output             i8_icb_rsp_err                ,
  output             i8_icb_rsp_excl_ok            ,
  output [  63:   0] i8_icb_rsp_rdata              ,
  output [   2:   0] i8_icb_rsp_usr                ,
    input              i9_icb_cmd_valid              ,
  output             i9_icb_cmd_ready              ,
  input              i9_icb_cmd_sel                ,
  input              i9_icb_cmd_read               ,
  input  [  31:   0] i9_icb_cmd_addr               ,
  input  [  63:   0] i9_icb_cmd_wdata              ,
  input  [   7:   0] i9_icb_cmd_wmask              ,
  input  [   2:   0] i9_icb_cmd_size               ,
  input              i9_icb_cmd_lock               ,
  input              i9_icb_cmd_excl               ,
  input  [   7:   0] i9_icb_cmd_xlen               ,
  input  [   1:   0] i9_icb_cmd_xburst             ,
  input  [   1:   0] i9_icb_cmd_modes              ,
  input              i9_icb_cmd_dmode              ,
  input  [   2:   0] i9_icb_cmd_attri              ,
  input  [   1:   0] i9_icb_cmd_beat               ,
  input  [   2:   0] i9_icb_cmd_usr                ,
  input              i9_icb_rsp_ready              ,
  output             i9_icb_rsp_valid              ,
  output             i9_icb_rsp_err                ,
  output             i9_icb_rsp_excl_ok            ,
  output [  63:   0] i9_icb_rsp_rdata              ,
  output [   2:   0] i9_icb_rsp_usr                ,
    input              i10_icb_cmd_valid             ,
  output             i10_icb_cmd_ready             ,
  input              i10_icb_cmd_sel               ,
  input              i10_icb_cmd_read              ,
  input  [  31:   0] i10_icb_cmd_addr              ,
  input  [  63:   0] i10_icb_cmd_wdata             ,
  input  [   7:   0] i10_icb_cmd_wmask             ,
  input  [   2:   0] i10_icb_cmd_size              ,
  input              i10_icb_cmd_lock              ,
  input              i10_icb_cmd_excl              ,
  input  [   7:   0] i10_icb_cmd_xlen              ,
  input  [   1:   0] i10_icb_cmd_xburst            ,
  input  [   1:   0] i10_icb_cmd_modes             ,
  input              i10_icb_cmd_dmode             ,
  input  [   2:   0] i10_icb_cmd_attri             ,
  input  [   1:   0] i10_icb_cmd_beat              ,
  input  [   2:   0] i10_icb_cmd_usr               ,
  input              i10_icb_rsp_ready             ,
  output             i10_icb_rsp_valid             ,
  output             i10_icb_rsp_err               ,
  output             i10_icb_rsp_excl_ok           ,
  output [  63:   0] i10_icb_rsp_rdata             ,
  output [   2:   0] i10_icb_rsp_usr               ,
    input              i11_icb_cmd_valid             ,
  output             i11_icb_cmd_ready             ,
  input              i11_icb_cmd_sel               ,
  input              i11_icb_cmd_read              ,
  input  [  31:   0] i11_icb_cmd_addr              ,
  input  [  63:   0] i11_icb_cmd_wdata             ,
  input  [   7:   0] i11_icb_cmd_wmask             ,
  input  [   2:   0] i11_icb_cmd_size              ,
  input              i11_icb_cmd_lock              ,
  input              i11_icb_cmd_excl              ,
  input  [   7:   0] i11_icb_cmd_xlen              ,
  input  [   1:   0] i11_icb_cmd_xburst            ,
  input  [   1:   0] i11_icb_cmd_modes             ,
  input              i11_icb_cmd_dmode             ,
  input  [   2:   0] i11_icb_cmd_attri             ,
  input  [   1:   0] i11_icb_cmd_beat              ,
  input  [   2:   0] i11_icb_cmd_usr               ,
  input              i11_icb_rsp_ready             ,
  output             i11_icb_rsp_valid             ,
  output             i11_icb_rsp_err               ,
  output             i11_icb_rsp_excl_ok           ,
  output [  63:   0] i11_icb_rsp_rdata             ,
  output [   2:   0] i11_icb_rsp_usr               ,
  input  clk,
  input  rst_n
  );
    wire    [  11:   0] arbt_bus_icb_cmd_valid        ;
  wire    [  11:   0] arbt_bus_icb_cmd_ready        ;
  wire    [  11:   0] arbt_bus_icb_cmd_sel          ;
  wire    [  11:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 767:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  95:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  35:   0] arbt_bus_icb_cmd_size         ;
  wire    [  11:   0] arbt_bus_icb_cmd_lock         ;
  wire    [  11:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  95:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  23:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  23:   0] arbt_bus_icb_cmd_modes        ;
  wire    [  11:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  35:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  23:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  35:   0] arbt_bus_icb_cmd_usr          ;
  wire    [  11:   0] arbt_bus_icb_rsp_ready        ;
  wire    [  11:   0] arbt_bus_icb_rsp_valid        ;
  wire    [  11:   0] arbt_bus_icb_rsp_err          ;
  wire    [  11:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 767:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  35:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i11_icb_cmd_valid
                           , i10_icb_cmd_valid
                           , i9_icb_cmd_valid
                           , i8_icb_cmd_valid
                           , i7_icb_cmd_valid
                           , i6_icb_cmd_valid
                           , i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i11_icb_cmd_sel
                           , i10_icb_cmd_sel
                           , i9_icb_cmd_sel
                           , i8_icb_cmd_sel
                           , i7_icb_cmd_sel
                           , i6_icb_cmd_sel
                           , i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i11_icb_cmd_read
                           , i10_icb_cmd_read
                           , i9_icb_cmd_read
                           , i8_icb_cmd_read
                           , i7_icb_cmd_read
                           , i6_icb_cmd_read
                           , i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i11_icb_cmd_addr
                           , i10_icb_cmd_addr
                           , i9_icb_cmd_addr
                           , i8_icb_cmd_addr
                           , i7_icb_cmd_addr
                           , i6_icb_cmd_addr
                           , i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i11_icb_cmd_wdata
                           , i10_icb_cmd_wdata
                           , i9_icb_cmd_wdata
                           , i8_icb_cmd_wdata
                           , i7_icb_cmd_wdata
                           , i6_icb_cmd_wdata
                           , i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i11_icb_cmd_wmask
                           , i10_icb_cmd_wmask
                           , i9_icb_cmd_wmask
                           , i8_icb_cmd_wmask
                           , i7_icb_cmd_wmask
                           , i6_icb_cmd_wmask
                           , i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i11_icb_cmd_size
                           , i10_icb_cmd_size
                           , i9_icb_cmd_size
                           , i8_icb_cmd_size
                           , i7_icb_cmd_size
                           , i6_icb_cmd_size
                           , i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i11_icb_cmd_lock
                           , i10_icb_cmd_lock
                           , i9_icb_cmd_lock
                           , i8_icb_cmd_lock
                           , i7_icb_cmd_lock
                           , i6_icb_cmd_lock
                           , i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i11_icb_cmd_excl
                           , i10_icb_cmd_excl
                           , i9_icb_cmd_excl
                           , i8_icb_cmd_excl
                           , i7_icb_cmd_excl
                           , i6_icb_cmd_excl
                           , i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i11_icb_cmd_xlen
                           , i10_icb_cmd_xlen
                           , i9_icb_cmd_xlen
                           , i8_icb_cmd_xlen
                           , i7_icb_cmd_xlen
                           , i6_icb_cmd_xlen
                           , i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i11_icb_cmd_xburst
                           , i10_icb_cmd_xburst
                           , i9_icb_cmd_xburst
                           , i8_icb_cmd_xburst
                           , i7_icb_cmd_xburst
                           , i6_icb_cmd_xburst
                           , i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i11_icb_cmd_modes
                           , i10_icb_cmd_modes
                           , i9_icb_cmd_modes
                           , i8_icb_cmd_modes
                           , i7_icb_cmd_modes
                           , i6_icb_cmd_modes
                           , i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i11_icb_cmd_dmode
                           , i10_icb_cmd_dmode
                           , i9_icb_cmd_dmode
                           , i8_icb_cmd_dmode
                           , i7_icb_cmd_dmode
                           , i6_icb_cmd_dmode
                           , i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i11_icb_cmd_attri
                           , i10_icb_cmd_attri
                           , i9_icb_cmd_attri
                           , i8_icb_cmd_attri
                           , i7_icb_cmd_attri
                           , i6_icb_cmd_attri
                           , i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i11_icb_cmd_beat
                           , i10_icb_cmd_beat
                           , i9_icb_cmd_beat
                           , i8_icb_cmd_beat
                           , i7_icb_cmd_beat
                           , i6_icb_cmd_beat
                           , i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i11_icb_cmd_usr
                           , i10_icb_cmd_usr
                           , i9_icb_cmd_usr
                           , i8_icb_cmd_usr
                           , i7_icb_cmd_usr
                           , i6_icb_cmd_usr
                           , i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i11_icb_cmd_ready
                           , i10_icb_cmd_ready
                           , i9_icb_cmd_ready
                           , i8_icb_cmd_ready
                           , i7_icb_cmd_ready
                           , i6_icb_cmd_ready
                           , i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i11_icb_rsp_valid
                           , i10_icb_rsp_valid
                           , i9_icb_rsp_valid
                           , i8_icb_rsp_valid
                           , i7_icb_rsp_valid
                           , i6_icb_rsp_valid
                           , i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i11_icb_rsp_err
                           , i10_icb_rsp_err
                           , i9_icb_rsp_err
                           , i8_icb_rsp_err
                           , i7_icb_rsp_err
                           , i6_icb_rsp_err
                           , i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i11_icb_rsp_excl_ok
                           , i10_icb_rsp_excl_ok
                           , i9_icb_rsp_excl_ok
                           , i8_icb_rsp_excl_ok
                           , i7_icb_rsp_excl_ok
                           , i6_icb_rsp_excl_ok
                           , i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i11_icb_rsp_rdata
                           , i10_icb_rsp_rdata
                           , i9_icb_rsp_rdata
                           , i8_icb_rsp_rdata
                           , i7_icb_rsp_rdata
                           , i6_icb_rsp_rdata
                           , i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i11_icb_rsp_usr
                           , i10_icb_rsp_usr
                           , i9_icb_rsp_usr
                           , i8_icb_rsp_usr
                           , i7_icb_rsp_usr
                           , i6_icb_rsp_usr
                           , i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i11_icb_rsp_ready
                           , i10_icb_rsp_ready
                           , i9_icb_rsp_ready
                           , i8_icb_rsp_ready
                           , i7_icb_rsp_ready
                           , i6_icb_rsp_ready
                           , i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (12),
  .ARBT_PTR_W (4),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [  11:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [  11:   0]),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read         [  11:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 383:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 767:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  95:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  35:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [  11:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [  11:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  95:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  23:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  23:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [  11:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  35:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  23:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  35:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [  11:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [  11:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [  11:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [  11:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 767:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  35:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv5_rw_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
    input              i6_icb_cmd_valid              ,
  output             i6_icb_cmd_ready              ,
  input              i6_icb_cmd_sel                ,
  input              i6_icb_cmd_read               ,
  input  [  31:   0] i6_icb_cmd_addr               ,
  input  [  63:   0] i6_icb_cmd_wdata              ,
  input  [   7:   0] i6_icb_cmd_wmask              ,
  input  [   2:   0] i6_icb_cmd_size               ,
  input              i6_icb_cmd_lock               ,
  input              i6_icb_cmd_excl               ,
  input  [   7:   0] i6_icb_cmd_xlen               ,
  input  [   1:   0] i6_icb_cmd_xburst             ,
  input  [   1:   0] i6_icb_cmd_modes              ,
  input              i6_icb_cmd_dmode              ,
  input  [   2:   0] i6_icb_cmd_attri              ,
  input  [   1:   0] i6_icb_cmd_beat               ,
  input  [   2:   0] i6_icb_cmd_usr                ,
  input              i6_icb_rsp_ready              ,
  output             i6_icb_rsp_valid              ,
  output             i6_icb_rsp_err                ,
  output             i6_icb_rsp_excl_ok            ,
  output [  63:   0] i6_icb_rsp_rdata              ,
  output [   2:   0] i6_icb_rsp_usr                ,
    input              i7_icb_cmd_valid              ,
  output             i7_icb_cmd_ready              ,
  input              i7_icb_cmd_sel                ,
  input              i7_icb_cmd_read               ,
  input  [  31:   0] i7_icb_cmd_addr               ,
  input  [  63:   0] i7_icb_cmd_wdata              ,
  input  [   7:   0] i7_icb_cmd_wmask              ,
  input  [   2:   0] i7_icb_cmd_size               ,
  input              i7_icb_cmd_lock               ,
  input              i7_icb_cmd_excl               ,
  input  [   7:   0] i7_icb_cmd_xlen               ,
  input  [   1:   0] i7_icb_cmd_xburst             ,
  input  [   1:   0] i7_icb_cmd_modes              ,
  input              i7_icb_cmd_dmode              ,
  input  [   2:   0] i7_icb_cmd_attri              ,
  input  [   1:   0] i7_icb_cmd_beat               ,
  input  [   2:   0] i7_icb_cmd_usr                ,
  input              i7_icb_rsp_ready              ,
  output             i7_icb_rsp_valid              ,
  output             i7_icb_rsp_err                ,
  output             i7_icb_rsp_excl_ok            ,
  output [  63:   0] i7_icb_rsp_rdata              ,
  output [   2:   0] i7_icb_rsp_usr                ,
    input              i8_icb_cmd_valid              ,
  output             i8_icb_cmd_ready              ,
  input              i8_icb_cmd_sel                ,
  input              i8_icb_cmd_read               ,
  input  [  31:   0] i8_icb_cmd_addr               ,
  input  [  63:   0] i8_icb_cmd_wdata              ,
  input  [   7:   0] i8_icb_cmd_wmask              ,
  input  [   2:   0] i8_icb_cmd_size               ,
  input              i8_icb_cmd_lock               ,
  input              i8_icb_cmd_excl               ,
  input  [   7:   0] i8_icb_cmd_xlen               ,
  input  [   1:   0] i8_icb_cmd_xburst             ,
  input  [   1:   0] i8_icb_cmd_modes              ,
  input              i8_icb_cmd_dmode              ,
  input  [   2:   0] i8_icb_cmd_attri              ,
  input  [   1:   0] i8_icb_cmd_beat               ,
  input  [   2:   0] i8_icb_cmd_usr                ,
  input              i8_icb_rsp_ready              ,
  output             i8_icb_rsp_valid              ,
  output             i8_icb_rsp_err                ,
  output             i8_icb_rsp_excl_ok            ,
  output [  63:   0] i8_icb_rsp_rdata              ,
  output [   2:   0] i8_icb_rsp_usr                ,
    input              i9_icb_cmd_valid              ,
  output             i9_icb_cmd_ready              ,
  input              i9_icb_cmd_sel                ,
  input              i9_icb_cmd_read               ,
  input  [  31:   0] i9_icb_cmd_addr               ,
  input  [  63:   0] i9_icb_cmd_wdata              ,
  input  [   7:   0] i9_icb_cmd_wmask              ,
  input  [   2:   0] i9_icb_cmd_size               ,
  input              i9_icb_cmd_lock               ,
  input              i9_icb_cmd_excl               ,
  input  [   7:   0] i9_icb_cmd_xlen               ,
  input  [   1:   0] i9_icb_cmd_xburst             ,
  input  [   1:   0] i9_icb_cmd_modes              ,
  input              i9_icb_cmd_dmode              ,
  input  [   2:   0] i9_icb_cmd_attri              ,
  input  [   1:   0] i9_icb_cmd_beat               ,
  input  [   2:   0] i9_icb_cmd_usr                ,
  input              i9_icb_rsp_ready              ,
  output             i9_icb_rsp_valid              ,
  output             i9_icb_rsp_err                ,
  output             i9_icb_rsp_excl_ok            ,
  output [  63:   0] i9_icb_rsp_rdata              ,
  output [   2:   0] i9_icb_rsp_usr                ,
    input              i10_icb_cmd_valid             ,
  output             i10_icb_cmd_ready             ,
  input              i10_icb_cmd_sel               ,
  input              i10_icb_cmd_read              ,
  input  [  31:   0] i10_icb_cmd_addr              ,
  input  [  63:   0] i10_icb_cmd_wdata             ,
  input  [   7:   0] i10_icb_cmd_wmask             ,
  input  [   2:   0] i10_icb_cmd_size              ,
  input              i10_icb_cmd_lock              ,
  input              i10_icb_cmd_excl              ,
  input  [   7:   0] i10_icb_cmd_xlen              ,
  input  [   1:   0] i10_icb_cmd_xburst            ,
  input  [   1:   0] i10_icb_cmd_modes             ,
  input              i10_icb_cmd_dmode             ,
  input  [   2:   0] i10_icb_cmd_attri             ,
  input  [   1:   0] i10_icb_cmd_beat              ,
  input  [   2:   0] i10_icb_cmd_usr               ,
  input              i10_icb_rsp_ready             ,
  output             i10_icb_rsp_valid             ,
  output             i10_icb_rsp_err               ,
  output             i10_icb_rsp_excl_ok           ,
  output [  63:   0] i10_icb_rsp_rdata             ,
  output [   2:   0] i10_icb_rsp_usr               ,
    input              i11_icb_cmd_valid             ,
  output             i11_icb_cmd_ready             ,
  input              i11_icb_cmd_sel               ,
  input              i11_icb_cmd_read              ,
  input  [  31:   0] i11_icb_cmd_addr              ,
  input  [  63:   0] i11_icb_cmd_wdata             ,
  input  [   7:   0] i11_icb_cmd_wmask             ,
  input  [   2:   0] i11_icb_cmd_size              ,
  input              i11_icb_cmd_lock              ,
  input              i11_icb_cmd_excl              ,
  input  [   7:   0] i11_icb_cmd_xlen              ,
  input  [   1:   0] i11_icb_cmd_xburst            ,
  input  [   1:   0] i11_icb_cmd_modes             ,
  input              i11_icb_cmd_dmode             ,
  input  [   2:   0] i11_icb_cmd_attri             ,
  input  [   1:   0] i11_icb_cmd_beat              ,
  input  [   2:   0] i11_icb_cmd_usr               ,
  input              i11_icb_rsp_ready             ,
  output             i11_icb_rsp_valid             ,
  output             i11_icb_rsp_err               ,
  output             i11_icb_rsp_excl_ok           ,
  output [  63:   0] i11_icb_rsp_rdata             ,
  output [   2:   0] i11_icb_rsp_usr               ,
  input  clk,
  input  rst_n
  );
    wire    [  11:   0] arbt_bus_icb_cmd_valid        ;
  wire    [  11:   0] arbt_bus_icb_cmd_ready        ;
  wire    [  11:   0] arbt_bus_icb_cmd_sel          ;
  wire    [  11:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 767:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  95:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  35:   0] arbt_bus_icb_cmd_size         ;
  wire    [  11:   0] arbt_bus_icb_cmd_lock         ;
  wire    [  11:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  95:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  23:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  23:   0] arbt_bus_icb_cmd_modes        ;
  wire    [  11:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  35:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  23:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  35:   0] arbt_bus_icb_cmd_usr          ;
  wire    [  11:   0] arbt_bus_icb_rsp_ready        ;
  wire    [  11:   0] arbt_bus_icb_rsp_valid        ;
  wire    [  11:   0] arbt_bus_icb_rsp_err          ;
  wire    [  11:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 767:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  35:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i11_icb_cmd_valid
                           , i10_icb_cmd_valid
                           , i9_icb_cmd_valid
                           , i8_icb_cmd_valid
                           , i7_icb_cmd_valid
                           , i6_icb_cmd_valid
                           , i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i11_icb_cmd_sel
                           , i10_icb_cmd_sel
                           , i9_icb_cmd_sel
                           , i8_icb_cmd_sel
                           , i7_icb_cmd_sel
                           , i6_icb_cmd_sel
                           , i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i11_icb_cmd_read
                           , i10_icb_cmd_read
                           , i9_icb_cmd_read
                           , i8_icb_cmd_read
                           , i7_icb_cmd_read
                           , i6_icb_cmd_read
                           , i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i11_icb_cmd_addr
                           , i10_icb_cmd_addr
                           , i9_icb_cmd_addr
                           , i8_icb_cmd_addr
                           , i7_icb_cmd_addr
                           , i6_icb_cmd_addr
                           , i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i11_icb_cmd_wdata
                           , i10_icb_cmd_wdata
                           , i9_icb_cmd_wdata
                           , i8_icb_cmd_wdata
                           , i7_icb_cmd_wdata
                           , i6_icb_cmd_wdata
                           , i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i11_icb_cmd_wmask
                           , i10_icb_cmd_wmask
                           , i9_icb_cmd_wmask
                           , i8_icb_cmd_wmask
                           , i7_icb_cmd_wmask
                           , i6_icb_cmd_wmask
                           , i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i11_icb_cmd_size
                           , i10_icb_cmd_size
                           , i9_icb_cmd_size
                           , i8_icb_cmd_size
                           , i7_icb_cmd_size
                           , i6_icb_cmd_size
                           , i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i11_icb_cmd_lock
                           , i10_icb_cmd_lock
                           , i9_icb_cmd_lock
                           , i8_icb_cmd_lock
                           , i7_icb_cmd_lock
                           , i6_icb_cmd_lock
                           , i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i11_icb_cmd_excl
                           , i10_icb_cmd_excl
                           , i9_icb_cmd_excl
                           , i8_icb_cmd_excl
                           , i7_icb_cmd_excl
                           , i6_icb_cmd_excl
                           , i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i11_icb_cmd_xlen
                           , i10_icb_cmd_xlen
                           , i9_icb_cmd_xlen
                           , i8_icb_cmd_xlen
                           , i7_icb_cmd_xlen
                           , i6_icb_cmd_xlen
                           , i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i11_icb_cmd_xburst
                           , i10_icb_cmd_xburst
                           , i9_icb_cmd_xburst
                           , i8_icb_cmd_xburst
                           , i7_icb_cmd_xburst
                           , i6_icb_cmd_xburst
                           , i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i11_icb_cmd_modes
                           , i10_icb_cmd_modes
                           , i9_icb_cmd_modes
                           , i8_icb_cmd_modes
                           , i7_icb_cmd_modes
                           , i6_icb_cmd_modes
                           , i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i11_icb_cmd_dmode
                           , i10_icb_cmd_dmode
                           , i9_icb_cmd_dmode
                           , i8_icb_cmd_dmode
                           , i7_icb_cmd_dmode
                           , i6_icb_cmd_dmode
                           , i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i11_icb_cmd_attri
                           , i10_icb_cmd_attri
                           , i9_icb_cmd_attri
                           , i8_icb_cmd_attri
                           , i7_icb_cmd_attri
                           , i6_icb_cmd_attri
                           , i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i11_icb_cmd_beat
                           , i10_icb_cmd_beat
                           , i9_icb_cmd_beat
                           , i8_icb_cmd_beat
                           , i7_icb_cmd_beat
                           , i6_icb_cmd_beat
                           , i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i11_icb_cmd_usr
                           , i10_icb_cmd_usr
                           , i9_icb_cmd_usr
                           , i8_icb_cmd_usr
                           , i7_icb_cmd_usr
                           , i6_icb_cmd_usr
                           , i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i11_icb_cmd_ready
                           , i10_icb_cmd_ready
                           , i9_icb_cmd_ready
                           , i8_icb_cmd_ready
                           , i7_icb_cmd_ready
                           , i6_icb_cmd_ready
                           , i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i11_icb_rsp_valid
                           , i10_icb_rsp_valid
                           , i9_icb_rsp_valid
                           , i8_icb_rsp_valid
                           , i7_icb_rsp_valid
                           , i6_icb_rsp_valid
                           , i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i11_icb_rsp_err
                           , i10_icb_rsp_err
                           , i9_icb_rsp_err
                           , i8_icb_rsp_err
                           , i7_icb_rsp_err
                           , i6_icb_rsp_err
                           , i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i11_icb_rsp_excl_ok
                           , i10_icb_rsp_excl_ok
                           , i9_icb_rsp_excl_ok
                           , i8_icb_rsp_excl_ok
                           , i7_icb_rsp_excl_ok
                           , i6_icb_rsp_excl_ok
                           , i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i11_icb_rsp_rdata
                           , i10_icb_rsp_rdata
                           , i9_icb_rsp_rdata
                           , i8_icb_rsp_rdata
                           , i7_icb_rsp_rdata
                           , i6_icb_rsp_rdata
                           , i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i11_icb_rsp_usr
                           , i10_icb_rsp_usr
                           , i9_icb_rsp_usr
                           , i8_icb_rsp_usr
                           , i7_icb_rsp_usr
                           , i6_icb_rsp_usr
                           , i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i11_icb_rsp_ready
                           , i10_icb_rsp_ready
                           , i9_icb_rsp_ready
                           , i8_icb_rsp_ready
                           , i7_icb_rsp_ready
                           , i6_icb_rsp_ready
                           , i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (12),
  .ARBT_PTR_W (4),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [  11:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [  11:   0]),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read         [  11:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 383:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 767:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  95:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  35:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [  11:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [  11:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  95:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  23:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  23:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [  11:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  35:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  23:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  35:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [  11:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [  11:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [  11:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [  11:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 767:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  35:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_xbar_slv6_rw_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
    input              i1_icb_cmd_valid              ,
  output             i1_icb_cmd_ready              ,
  input              i1_icb_cmd_sel                ,
  input              i1_icb_cmd_read               ,
  input  [  31:   0] i1_icb_cmd_addr               ,
  input  [  63:   0] i1_icb_cmd_wdata              ,
  input  [   7:   0] i1_icb_cmd_wmask              ,
  input  [   2:   0] i1_icb_cmd_size               ,
  input              i1_icb_cmd_lock               ,
  input              i1_icb_cmd_excl               ,
  input  [   7:   0] i1_icb_cmd_xlen               ,
  input  [   1:   0] i1_icb_cmd_xburst             ,
  input  [   1:   0] i1_icb_cmd_modes              ,
  input              i1_icb_cmd_dmode              ,
  input  [   2:   0] i1_icb_cmd_attri              ,
  input  [   1:   0] i1_icb_cmd_beat               ,
  input  [   2:   0] i1_icb_cmd_usr                ,
  input              i1_icb_rsp_ready              ,
  output             i1_icb_rsp_valid              ,
  output             i1_icb_rsp_err                ,
  output             i1_icb_rsp_excl_ok            ,
  output [  63:   0] i1_icb_rsp_rdata              ,
  output [   2:   0] i1_icb_rsp_usr                ,
    input              i2_icb_cmd_valid              ,
  output             i2_icb_cmd_ready              ,
  input              i2_icb_cmd_sel                ,
  input              i2_icb_cmd_read               ,
  input  [  31:   0] i2_icb_cmd_addr               ,
  input  [  63:   0] i2_icb_cmd_wdata              ,
  input  [   7:   0] i2_icb_cmd_wmask              ,
  input  [   2:   0] i2_icb_cmd_size               ,
  input              i2_icb_cmd_lock               ,
  input              i2_icb_cmd_excl               ,
  input  [   7:   0] i2_icb_cmd_xlen               ,
  input  [   1:   0] i2_icb_cmd_xburst             ,
  input  [   1:   0] i2_icb_cmd_modes              ,
  input              i2_icb_cmd_dmode              ,
  input  [   2:   0] i2_icb_cmd_attri              ,
  input  [   1:   0] i2_icb_cmd_beat               ,
  input  [   2:   0] i2_icb_cmd_usr                ,
  input              i2_icb_rsp_ready              ,
  output             i2_icb_rsp_valid              ,
  output             i2_icb_rsp_err                ,
  output             i2_icb_rsp_excl_ok            ,
  output [  63:   0] i2_icb_rsp_rdata              ,
  output [   2:   0] i2_icb_rsp_usr                ,
    input              i3_icb_cmd_valid              ,
  output             i3_icb_cmd_ready              ,
  input              i3_icb_cmd_sel                ,
  input              i3_icb_cmd_read               ,
  input  [  31:   0] i3_icb_cmd_addr               ,
  input  [  63:   0] i3_icb_cmd_wdata              ,
  input  [   7:   0] i3_icb_cmd_wmask              ,
  input  [   2:   0] i3_icb_cmd_size               ,
  input              i3_icb_cmd_lock               ,
  input              i3_icb_cmd_excl               ,
  input  [   7:   0] i3_icb_cmd_xlen               ,
  input  [   1:   0] i3_icb_cmd_xburst             ,
  input  [   1:   0] i3_icb_cmd_modes              ,
  input              i3_icb_cmd_dmode              ,
  input  [   2:   0] i3_icb_cmd_attri              ,
  input  [   1:   0] i3_icb_cmd_beat               ,
  input  [   2:   0] i3_icb_cmd_usr                ,
  input              i3_icb_rsp_ready              ,
  output             i3_icb_rsp_valid              ,
  output             i3_icb_rsp_err                ,
  output             i3_icb_rsp_excl_ok            ,
  output [  63:   0] i3_icb_rsp_rdata              ,
  output [   2:   0] i3_icb_rsp_usr                ,
    input              i4_icb_cmd_valid              ,
  output             i4_icb_cmd_ready              ,
  input              i4_icb_cmd_sel                ,
  input              i4_icb_cmd_read               ,
  input  [  31:   0] i4_icb_cmd_addr               ,
  input  [  63:   0] i4_icb_cmd_wdata              ,
  input  [   7:   0] i4_icb_cmd_wmask              ,
  input  [   2:   0] i4_icb_cmd_size               ,
  input              i4_icb_cmd_lock               ,
  input              i4_icb_cmd_excl               ,
  input  [   7:   0] i4_icb_cmd_xlen               ,
  input  [   1:   0] i4_icb_cmd_xburst             ,
  input  [   1:   0] i4_icb_cmd_modes              ,
  input              i4_icb_cmd_dmode              ,
  input  [   2:   0] i4_icb_cmd_attri              ,
  input  [   1:   0] i4_icb_cmd_beat               ,
  input  [   2:   0] i4_icb_cmd_usr                ,
  input              i4_icb_rsp_ready              ,
  output             i4_icb_rsp_valid              ,
  output             i4_icb_rsp_err                ,
  output             i4_icb_rsp_excl_ok            ,
  output [  63:   0] i4_icb_rsp_rdata              ,
  output [   2:   0] i4_icb_rsp_usr                ,
    input              i5_icb_cmd_valid              ,
  output             i5_icb_cmd_ready              ,
  input              i5_icb_cmd_sel                ,
  input              i5_icb_cmd_read               ,
  input  [  31:   0] i5_icb_cmd_addr               ,
  input  [  63:   0] i5_icb_cmd_wdata              ,
  input  [   7:   0] i5_icb_cmd_wmask              ,
  input  [   2:   0] i5_icb_cmd_size               ,
  input              i5_icb_cmd_lock               ,
  input              i5_icb_cmd_excl               ,
  input  [   7:   0] i5_icb_cmd_xlen               ,
  input  [   1:   0] i5_icb_cmd_xburst             ,
  input  [   1:   0] i5_icb_cmd_modes              ,
  input              i5_icb_cmd_dmode              ,
  input  [   2:   0] i5_icb_cmd_attri              ,
  input  [   1:   0] i5_icb_cmd_beat               ,
  input  [   2:   0] i5_icb_cmd_usr                ,
  input              i5_icb_rsp_ready              ,
  output             i5_icb_rsp_valid              ,
  output             i5_icb_rsp_err                ,
  output             i5_icb_rsp_excl_ok            ,
  output [  63:   0] i5_icb_rsp_rdata              ,
  output [   2:   0] i5_icb_rsp_usr                ,
    input              i6_icb_cmd_valid              ,
  output             i6_icb_cmd_ready              ,
  input              i6_icb_cmd_sel                ,
  input              i6_icb_cmd_read               ,
  input  [  31:   0] i6_icb_cmd_addr               ,
  input  [  63:   0] i6_icb_cmd_wdata              ,
  input  [   7:   0] i6_icb_cmd_wmask              ,
  input  [   2:   0] i6_icb_cmd_size               ,
  input              i6_icb_cmd_lock               ,
  input              i6_icb_cmd_excl               ,
  input  [   7:   0] i6_icb_cmd_xlen               ,
  input  [   1:   0] i6_icb_cmd_xburst             ,
  input  [   1:   0] i6_icb_cmd_modes              ,
  input              i6_icb_cmd_dmode              ,
  input  [   2:   0] i6_icb_cmd_attri              ,
  input  [   1:   0] i6_icb_cmd_beat               ,
  input  [   2:   0] i6_icb_cmd_usr                ,
  input              i6_icb_rsp_ready              ,
  output             i6_icb_rsp_valid              ,
  output             i6_icb_rsp_err                ,
  output             i6_icb_rsp_excl_ok            ,
  output [  63:   0] i6_icb_rsp_rdata              ,
  output [   2:   0] i6_icb_rsp_usr                ,
    input              i7_icb_cmd_valid              ,
  output             i7_icb_cmd_ready              ,
  input              i7_icb_cmd_sel                ,
  input              i7_icb_cmd_read               ,
  input  [  31:   0] i7_icb_cmd_addr               ,
  input  [  63:   0] i7_icb_cmd_wdata              ,
  input  [   7:   0] i7_icb_cmd_wmask              ,
  input  [   2:   0] i7_icb_cmd_size               ,
  input              i7_icb_cmd_lock               ,
  input              i7_icb_cmd_excl               ,
  input  [   7:   0] i7_icb_cmd_xlen               ,
  input  [   1:   0] i7_icb_cmd_xburst             ,
  input  [   1:   0] i7_icb_cmd_modes              ,
  input              i7_icb_cmd_dmode              ,
  input  [   2:   0] i7_icb_cmd_attri              ,
  input  [   1:   0] i7_icb_cmd_beat               ,
  input  [   2:   0] i7_icb_cmd_usr                ,
  input              i7_icb_rsp_ready              ,
  output             i7_icb_rsp_valid              ,
  output             i7_icb_rsp_err                ,
  output             i7_icb_rsp_excl_ok            ,
  output [  63:   0] i7_icb_rsp_rdata              ,
  output [   2:   0] i7_icb_rsp_usr                ,
    input              i8_icb_cmd_valid              ,
  output             i8_icb_cmd_ready              ,
  input              i8_icb_cmd_sel                ,
  input              i8_icb_cmd_read               ,
  input  [  31:   0] i8_icb_cmd_addr               ,
  input  [  63:   0] i8_icb_cmd_wdata              ,
  input  [   7:   0] i8_icb_cmd_wmask              ,
  input  [   2:   0] i8_icb_cmd_size               ,
  input              i8_icb_cmd_lock               ,
  input              i8_icb_cmd_excl               ,
  input  [   7:   0] i8_icb_cmd_xlen               ,
  input  [   1:   0] i8_icb_cmd_xburst             ,
  input  [   1:   0] i8_icb_cmd_modes              ,
  input              i8_icb_cmd_dmode              ,
  input  [   2:   0] i8_icb_cmd_attri              ,
  input  [   1:   0] i8_icb_cmd_beat               ,
  input  [   2:   0] i8_icb_cmd_usr                ,
  input              i8_icb_rsp_ready              ,
  output             i8_icb_rsp_valid              ,
  output             i8_icb_rsp_err                ,
  output             i8_icb_rsp_excl_ok            ,
  output [  63:   0] i8_icb_rsp_rdata              ,
  output [   2:   0] i8_icb_rsp_usr                ,
    input              i9_icb_cmd_valid              ,
  output             i9_icb_cmd_ready              ,
  input              i9_icb_cmd_sel                ,
  input              i9_icb_cmd_read               ,
  input  [  31:   0] i9_icb_cmd_addr               ,
  input  [  63:   0] i9_icb_cmd_wdata              ,
  input  [   7:   0] i9_icb_cmd_wmask              ,
  input  [   2:   0] i9_icb_cmd_size               ,
  input              i9_icb_cmd_lock               ,
  input              i9_icb_cmd_excl               ,
  input  [   7:   0] i9_icb_cmd_xlen               ,
  input  [   1:   0] i9_icb_cmd_xburst             ,
  input  [   1:   0] i9_icb_cmd_modes              ,
  input              i9_icb_cmd_dmode              ,
  input  [   2:   0] i9_icb_cmd_attri              ,
  input  [   1:   0] i9_icb_cmd_beat               ,
  input  [   2:   0] i9_icb_cmd_usr                ,
  input              i9_icb_rsp_ready              ,
  output             i9_icb_rsp_valid              ,
  output             i9_icb_rsp_err                ,
  output             i9_icb_rsp_excl_ok            ,
  output [  63:   0] i9_icb_rsp_rdata              ,
  output [   2:   0] i9_icb_rsp_usr                ,
    input              i10_icb_cmd_valid             ,
  output             i10_icb_cmd_ready             ,
  input              i10_icb_cmd_sel               ,
  input              i10_icb_cmd_read              ,
  input  [  31:   0] i10_icb_cmd_addr              ,
  input  [  63:   0] i10_icb_cmd_wdata             ,
  input  [   7:   0] i10_icb_cmd_wmask             ,
  input  [   2:   0] i10_icb_cmd_size              ,
  input              i10_icb_cmd_lock              ,
  input              i10_icb_cmd_excl              ,
  input  [   7:   0] i10_icb_cmd_xlen              ,
  input  [   1:   0] i10_icb_cmd_xburst            ,
  input  [   1:   0] i10_icb_cmd_modes             ,
  input              i10_icb_cmd_dmode             ,
  input  [   2:   0] i10_icb_cmd_attri             ,
  input  [   1:   0] i10_icb_cmd_beat              ,
  input  [   2:   0] i10_icb_cmd_usr               ,
  input              i10_icb_rsp_ready             ,
  output             i10_icb_rsp_valid             ,
  output             i10_icb_rsp_err               ,
  output             i10_icb_rsp_excl_ok           ,
  output [  63:   0] i10_icb_rsp_rdata             ,
  output [   2:   0] i10_icb_rsp_usr               ,
    input              i11_icb_cmd_valid             ,
  output             i11_icb_cmd_ready             ,
  input              i11_icb_cmd_sel               ,
  input              i11_icb_cmd_read              ,
  input  [  31:   0] i11_icb_cmd_addr              ,
  input  [  63:   0] i11_icb_cmd_wdata             ,
  input  [   7:   0] i11_icb_cmd_wmask             ,
  input  [   2:   0] i11_icb_cmd_size              ,
  input              i11_icb_cmd_lock              ,
  input              i11_icb_cmd_excl              ,
  input  [   7:   0] i11_icb_cmd_xlen              ,
  input  [   1:   0] i11_icb_cmd_xburst            ,
  input  [   1:   0] i11_icb_cmd_modes             ,
  input              i11_icb_cmd_dmode             ,
  input  [   2:   0] i11_icb_cmd_attri             ,
  input  [   1:   0] i11_icb_cmd_beat              ,
  input  [   2:   0] i11_icb_cmd_usr               ,
  input              i11_icb_rsp_ready             ,
  output             i11_icb_rsp_valid             ,
  output             i11_icb_rsp_err               ,
  output             i11_icb_rsp_excl_ok           ,
  output [  63:   0] i11_icb_rsp_rdata             ,
  output [   2:   0] i11_icb_rsp_usr               ,
  input  clk,
  input  rst_n
  );
    wire    [  11:   0] arbt_bus_icb_cmd_valid        ;
  wire    [  11:   0] arbt_bus_icb_cmd_ready        ;
  wire    [  11:   0] arbt_bus_icb_cmd_sel          ;
  wire    [  11:   0] arbt_bus_icb_cmd_read         ;
  wire    [ 383:   0] arbt_bus_icb_cmd_addr         ;
  wire    [ 767:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [  95:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [  35:   0] arbt_bus_icb_cmd_size         ;
  wire    [  11:   0] arbt_bus_icb_cmd_lock         ;
  wire    [  11:   0] arbt_bus_icb_cmd_excl         ;
  wire    [  95:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [  23:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [  23:   0] arbt_bus_icb_cmd_modes        ;
  wire    [  11:   0] arbt_bus_icb_cmd_dmode        ;
  wire    [  35:   0] arbt_bus_icb_cmd_attri        ;
  wire    [  23:   0] arbt_bus_icb_cmd_beat         ;
  wire    [  35:   0] arbt_bus_icb_cmd_usr          ;
  wire    [  11:   0] arbt_bus_icb_rsp_ready        ;
  wire    [  11:   0] arbt_bus_icb_rsp_valid        ;
  wire    [  11:   0] arbt_bus_icb_rsp_err          ;
  wire    [  11:   0] arbt_bus_icb_rsp_excl_ok      ;
  wire    [ 767:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [  35:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i11_icb_cmd_valid
                           , i10_icb_cmd_valid
                           , i9_icb_cmd_valid
                           , i8_icb_cmd_valid
                           , i7_icb_cmd_valid
                           , i6_icb_cmd_valid
                           , i5_icb_cmd_valid
                           , i4_icb_cmd_valid
                           , i3_icb_cmd_valid
                           , i2_icb_cmd_valid
                           , i1_icb_cmd_valid
                           , i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i11_icb_cmd_sel
                           , i10_icb_cmd_sel
                           , i9_icb_cmd_sel
                           , i8_icb_cmd_sel
                           , i7_icb_cmd_sel
                           , i6_icb_cmd_sel
                           , i5_icb_cmd_sel
                           , i4_icb_cmd_sel
                           , i3_icb_cmd_sel
                           , i2_icb_cmd_sel
                           , i1_icb_cmd_sel
                           , i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i11_icb_cmd_read
                           , i10_icb_cmd_read
                           , i9_icb_cmd_read
                           , i8_icb_cmd_read
                           , i7_icb_cmd_read
                           , i6_icb_cmd_read
                           , i5_icb_cmd_read
                           , i4_icb_cmd_read
                           , i3_icb_cmd_read
                           , i2_icb_cmd_read
                           , i1_icb_cmd_read
                           , i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i11_icb_cmd_addr
                           , i10_icb_cmd_addr
                           , i9_icb_cmd_addr
                           , i8_icb_cmd_addr
                           , i7_icb_cmd_addr
                           , i6_icb_cmd_addr
                           , i5_icb_cmd_addr
                           , i4_icb_cmd_addr
                           , i3_icb_cmd_addr
                           , i2_icb_cmd_addr
                           , i1_icb_cmd_addr
                           , i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i11_icb_cmd_wdata
                           , i10_icb_cmd_wdata
                           , i9_icb_cmd_wdata
                           , i8_icb_cmd_wdata
                           , i7_icb_cmd_wdata
                           , i6_icb_cmd_wdata
                           , i5_icb_cmd_wdata
                           , i4_icb_cmd_wdata
                           , i3_icb_cmd_wdata
                           , i2_icb_cmd_wdata
                           , i1_icb_cmd_wdata
                           , i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i11_icb_cmd_wmask
                           , i10_icb_cmd_wmask
                           , i9_icb_cmd_wmask
                           , i8_icb_cmd_wmask
                           , i7_icb_cmd_wmask
                           , i6_icb_cmd_wmask
                           , i5_icb_cmd_wmask
                           , i4_icb_cmd_wmask
                           , i3_icb_cmd_wmask
                           , i2_icb_cmd_wmask
                           , i1_icb_cmd_wmask
                           , i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i11_icb_cmd_size
                           , i10_icb_cmd_size
                           , i9_icb_cmd_size
                           , i8_icb_cmd_size
                           , i7_icb_cmd_size
                           , i6_icb_cmd_size
                           , i5_icb_cmd_size
                           , i4_icb_cmd_size
                           , i3_icb_cmd_size
                           , i2_icb_cmd_size
                           , i1_icb_cmd_size
                           , i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i11_icb_cmd_lock
                           , i10_icb_cmd_lock
                           , i9_icb_cmd_lock
                           , i8_icb_cmd_lock
                           , i7_icb_cmd_lock
                           , i6_icb_cmd_lock
                           , i5_icb_cmd_lock
                           , i4_icb_cmd_lock
                           , i3_icb_cmd_lock
                           , i2_icb_cmd_lock
                           , i1_icb_cmd_lock
                           , i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i11_icb_cmd_excl
                           , i10_icb_cmd_excl
                           , i9_icb_cmd_excl
                           , i8_icb_cmd_excl
                           , i7_icb_cmd_excl
                           , i6_icb_cmd_excl
                           , i5_icb_cmd_excl
                           , i4_icb_cmd_excl
                           , i3_icb_cmd_excl
                           , i2_icb_cmd_excl
                           , i1_icb_cmd_excl
                           , i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i11_icb_cmd_xlen
                           , i10_icb_cmd_xlen
                           , i9_icb_cmd_xlen
                           , i8_icb_cmd_xlen
                           , i7_icb_cmd_xlen
                           , i6_icb_cmd_xlen
                           , i5_icb_cmd_xlen
                           , i4_icb_cmd_xlen
                           , i3_icb_cmd_xlen
                           , i2_icb_cmd_xlen
                           , i1_icb_cmd_xlen
                           , i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i11_icb_cmd_xburst
                           , i10_icb_cmd_xburst
                           , i9_icb_cmd_xburst
                           , i8_icb_cmd_xburst
                           , i7_icb_cmd_xburst
                           , i6_icb_cmd_xburst
                           , i5_icb_cmd_xburst
                           , i4_icb_cmd_xburst
                           , i3_icb_cmd_xburst
                           , i2_icb_cmd_xburst
                           , i1_icb_cmd_xburst
                           , i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i11_icb_cmd_modes
                           , i10_icb_cmd_modes
                           , i9_icb_cmd_modes
                           , i8_icb_cmd_modes
                           , i7_icb_cmd_modes
                           , i6_icb_cmd_modes
                           , i5_icb_cmd_modes
                           , i4_icb_cmd_modes
                           , i3_icb_cmd_modes
                           , i2_icb_cmd_modes
                           , i1_icb_cmd_modes
                           , i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i11_icb_cmd_dmode
                           , i10_icb_cmd_dmode
                           , i9_icb_cmd_dmode
                           , i8_icb_cmd_dmode
                           , i7_icb_cmd_dmode
                           , i6_icb_cmd_dmode
                           , i5_icb_cmd_dmode
                           , i4_icb_cmd_dmode
                           , i3_icb_cmd_dmode
                           , i2_icb_cmd_dmode
                           , i1_icb_cmd_dmode
                           , i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i11_icb_cmd_attri
                           , i10_icb_cmd_attri
                           , i9_icb_cmd_attri
                           , i8_icb_cmd_attri
                           , i7_icb_cmd_attri
                           , i6_icb_cmd_attri
                           , i5_icb_cmd_attri
                           , i4_icb_cmd_attri
                           , i3_icb_cmd_attri
                           , i2_icb_cmd_attri
                           , i1_icb_cmd_attri
                           , i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i11_icb_cmd_beat
                           , i10_icb_cmd_beat
                           , i9_icb_cmd_beat
                           , i8_icb_cmd_beat
                           , i7_icb_cmd_beat
                           , i6_icb_cmd_beat
                           , i5_icb_cmd_beat
                           , i4_icb_cmd_beat
                           , i3_icb_cmd_beat
                           , i2_icb_cmd_beat
                           , i1_icb_cmd_beat
                           , i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i11_icb_cmd_usr
                           , i10_icb_cmd_usr
                           , i9_icb_cmd_usr
                           , i8_icb_cmd_usr
                           , i7_icb_cmd_usr
                           , i6_icb_cmd_usr
                           , i5_icb_cmd_usr
                           , i4_icb_cmd_usr
                           , i3_icb_cmd_usr
                           , i2_icb_cmd_usr
                           , i1_icb_cmd_usr
                           , i0_icb_cmd_usr
                           };
      assign                 { i11_icb_cmd_ready
                           , i10_icb_cmd_ready
                           , i9_icb_cmd_ready
                           , i8_icb_cmd_ready
                           , i7_icb_cmd_ready
                           , i6_icb_cmd_ready
                           , i5_icb_cmd_ready
                           , i4_icb_cmd_ready
                           , i3_icb_cmd_ready
                           , i2_icb_cmd_ready
                           , i1_icb_cmd_ready
                           , i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i11_icb_rsp_valid
                           , i10_icb_rsp_valid
                           , i9_icb_rsp_valid
                           , i8_icb_rsp_valid
                           , i7_icb_rsp_valid
                           , i6_icb_rsp_valid
                           , i5_icb_rsp_valid
                           , i4_icb_rsp_valid
                           , i3_icb_rsp_valid
                           , i2_icb_rsp_valid
                           , i1_icb_rsp_valid
                           , i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i11_icb_rsp_err
                           , i10_icb_rsp_err
                           , i9_icb_rsp_err
                           , i8_icb_rsp_err
                           , i7_icb_rsp_err
                           , i6_icb_rsp_err
                           , i5_icb_rsp_err
                           , i4_icb_rsp_err
                           , i3_icb_rsp_err
                           , i2_icb_rsp_err
                           , i1_icb_rsp_err
                           , i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i11_icb_rsp_excl_ok
                           , i10_icb_rsp_excl_ok
                           , i9_icb_rsp_excl_ok
                           , i8_icb_rsp_excl_ok
                           , i7_icb_rsp_excl_ok
                           , i6_icb_rsp_excl_ok
                           , i5_icb_rsp_excl_ok
                           , i4_icb_rsp_excl_ok
                           , i3_icb_rsp_excl_ok
                           , i2_icb_rsp_excl_ok
                           , i1_icb_rsp_excl_ok
                           , i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i11_icb_rsp_rdata
                           , i10_icb_rsp_rdata
                           , i9_icb_rsp_rdata
                           , i8_icb_rsp_rdata
                           , i7_icb_rsp_rdata
                           , i6_icb_rsp_rdata
                           , i5_icb_rsp_rdata
                           , i4_icb_rsp_rdata
                           , i3_icb_rsp_rdata
                           , i2_icb_rsp_rdata
                           , i1_icb_rsp_rdata
                           , i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i11_icb_rsp_usr
                           , i10_icb_rsp_usr
                           , i9_icb_rsp_usr
                           , i8_icb_rsp_usr
                           , i7_icb_rsp_usr
                           , i6_icb_rsp_usr
                           , i5_icb_rsp_usr
                           , i4_icb_rsp_usr
                           , i3_icb_rsp_usr
                           , i2_icb_rsp_usr
                           , i1_icb_rsp_usr
                           , i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i11_icb_rsp_ready
                           , i10_icb_rsp_ready
                           , i9_icb_rsp_ready
                           , i8_icb_rsp_ready
                           , i7_icb_rsp_ready
                           , i6_icb_rsp_ready
                           , i5_icb_rsp_ready
                           , i4_icb_rsp_ready
                           , i3_icb_rsp_ready
                           , i2_icb_rsp_ready
                           , i1_icb_rsp_ready
                           , i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (12),
  .ARBT_PTR_W (4),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid        [  11:   0]),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready        [  11:   0]),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read         [  11:   0]),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [ 383:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [ 767:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [  95:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [  35:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock         [  11:   0]),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl         [  11:   0]),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [  95:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [  23:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [  23:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode        [  11:   0]),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [  35:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [  23:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [  35:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready        [  11:   0]),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid        [  11:   0]),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err          [  11:   0]),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok      [  11:   0]),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [ 767:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [  35:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_mgrp0_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                arbt_bus_icb_cmd_valid        ;
  wire                arbt_bus_icb_cmd_ready        ;
  wire                arbt_bus_icb_cmd_sel          ;
  wire                arbt_bus_icb_cmd_read         ;
  wire    [  31:   0] arbt_bus_icb_cmd_addr         ;
  wire    [  63:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] arbt_bus_icb_cmd_size         ;
  wire                arbt_bus_icb_cmd_lock         ;
  wire                arbt_bus_icb_cmd_excl         ;
  wire    [   7:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] arbt_bus_icb_cmd_modes        ;
  wire                arbt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] arbt_bus_icb_cmd_attri        ;
  wire    [   1:   0] arbt_bus_icb_cmd_beat         ;
  wire    [   2:   0] arbt_bus_icb_cmd_usr          ;
  wire                arbt_bus_icb_rsp_ready        ;
  wire                arbt_bus_icb_rsp_valid        ;
  wire                arbt_bus_icb_rsp_err          ;
  wire                arbt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i0_icb_cmd_usr
                           };
      assign                 { i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (1),
  .ARBT_PTR_W (1),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid                   ),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready                   ),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read                    ),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [  31:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [  63:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [   7:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [   2:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock                    ),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl                    ),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [   7:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [   1:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [   1:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode                   ),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [   2:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [   1:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [   2:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready                   ),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid                   ),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err                     ),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok                 ),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [  63:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [   2:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_mgrp1_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                arbt_bus_icb_cmd_valid        ;
  wire                arbt_bus_icb_cmd_ready        ;
  wire                arbt_bus_icb_cmd_sel          ;
  wire                arbt_bus_icb_cmd_read         ;
  wire    [  31:   0] arbt_bus_icb_cmd_addr         ;
  wire    [  63:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] arbt_bus_icb_cmd_size         ;
  wire                arbt_bus_icb_cmd_lock         ;
  wire                arbt_bus_icb_cmd_excl         ;
  wire    [   7:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] arbt_bus_icb_cmd_modes        ;
  wire                arbt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] arbt_bus_icb_cmd_attri        ;
  wire    [   1:   0] arbt_bus_icb_cmd_beat         ;
  wire    [   2:   0] arbt_bus_icb_cmd_usr          ;
  wire                arbt_bus_icb_rsp_ready        ;
  wire                arbt_bus_icb_rsp_valid        ;
  wire                arbt_bus_icb_rsp_err          ;
  wire                arbt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i0_icb_cmd_usr
                           };
      assign                 { i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (1),
  .ARBT_PTR_W (1),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_read (1'b1),
    .i_bus_icb_cmd_wdata({(64*1){1'b0}}),
    .i_bus_icb_cmd_wmask({((64*1)/8){1'b0}}),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid                   ),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready                   ),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [  31:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [   2:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock                    ),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl                    ),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [   7:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [   1:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [   1:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode                   ),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [   2:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [   1:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [   2:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready                   ),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid                   ),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err                     ),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok                 ),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [  63:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [   2:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_read (1'b1),
    .i_icb_cmd_wdata(64'b0),
    .i_icb_cmd_wmask({64/8{1'b0}}),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_mgrp2_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                arbt_bus_icb_cmd_valid        ;
  wire                arbt_bus_icb_cmd_ready        ;
  wire                arbt_bus_icb_cmd_sel          ;
  wire                arbt_bus_icb_cmd_read         ;
  wire    [  31:   0] arbt_bus_icb_cmd_addr         ;
  wire    [  63:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] arbt_bus_icb_cmd_size         ;
  wire                arbt_bus_icb_cmd_lock         ;
  wire                arbt_bus_icb_cmd_excl         ;
  wire    [   7:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] arbt_bus_icb_cmd_modes        ;
  wire                arbt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] arbt_bus_icb_cmd_attri        ;
  wire    [   1:   0] arbt_bus_icb_cmd_beat         ;
  wire    [   2:   0] arbt_bus_icb_cmd_usr          ;
  wire                arbt_bus_icb_rsp_ready        ;
  wire                arbt_bus_icb_rsp_valid        ;
  wire                arbt_bus_icb_rsp_err          ;
  wire                arbt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i0_icb_cmd_usr
                           };
      assign                 { i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (1),
  .ARBT_PTR_W (1),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
    .i_bus_icb_cmd_read (1'b0),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid                   ),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready                   ),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [  31:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [  63:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [   7:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [   2:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock                    ),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl                    ),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [   7:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [   1:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [   1:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode                   ),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [   2:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [   1:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [   2:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready                   ),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid                   ),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err                     ),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok                 ),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [  63:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
    .i_icb_cmd_read (1'b0),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .o_icb_rsp_rdata(64'b0),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_mgrp3_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                arbt_bus_icb_cmd_valid        ;
  wire                arbt_bus_icb_cmd_ready        ;
  wire                arbt_bus_icb_cmd_sel          ;
  wire                arbt_bus_icb_cmd_read         ;
  wire    [  31:   0] arbt_bus_icb_cmd_addr         ;
  wire    [  63:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] arbt_bus_icb_cmd_size         ;
  wire                arbt_bus_icb_cmd_lock         ;
  wire                arbt_bus_icb_cmd_excl         ;
  wire    [   7:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] arbt_bus_icb_cmd_modes        ;
  wire                arbt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] arbt_bus_icb_cmd_attri        ;
  wire    [   1:   0] arbt_bus_icb_cmd_beat         ;
  wire    [   2:   0] arbt_bus_icb_cmd_usr          ;
  wire                arbt_bus_icb_rsp_ready        ;
  wire                arbt_bus_icb_rsp_valid        ;
  wire                arbt_bus_icb_rsp_err          ;
  wire                arbt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i0_icb_cmd_usr
                           };
      assign                 { i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (1),
  .ARBT_PTR_W (1),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid                   ),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready                   ),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read                    ),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [  31:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [  63:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [   7:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [   2:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock                    ),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl                    ),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [   7:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [   1:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [   1:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode                   ),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [   2:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [   1:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [   2:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready                   ),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid                   ),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err                     ),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok                 ),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [  63:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [   2:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_mgrp4_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                arbt_bus_icb_cmd_valid        ;
  wire                arbt_bus_icb_cmd_ready        ;
  wire                arbt_bus_icb_cmd_sel          ;
  wire                arbt_bus_icb_cmd_read         ;
  wire    [  31:   0] arbt_bus_icb_cmd_addr         ;
  wire    [  63:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] arbt_bus_icb_cmd_size         ;
  wire                arbt_bus_icb_cmd_lock         ;
  wire                arbt_bus_icb_cmd_excl         ;
  wire    [   7:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] arbt_bus_icb_cmd_modes        ;
  wire                arbt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] arbt_bus_icb_cmd_attri        ;
  wire    [   1:   0] arbt_bus_icb_cmd_beat         ;
  wire    [   2:   0] arbt_bus_icb_cmd_usr          ;
  wire                arbt_bus_icb_rsp_ready        ;
  wire                arbt_bus_icb_rsp_valid        ;
  wire                arbt_bus_icb_rsp_err          ;
  wire                arbt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i0_icb_cmd_usr
                           };
      assign                 { i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (1),
  .ARBT_PTR_W (1),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid                   ),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready                   ),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read                    ),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [  31:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [  63:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [   7:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [   2:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock                    ),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl                    ),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [   7:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [   1:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [   1:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode                   ),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [   2:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [   1:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [   2:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready                   ),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid                   ),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err                     ),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok                 ),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [  63:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [   2:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_mgrp5_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                arbt_bus_icb_cmd_valid        ;
  wire                arbt_bus_icb_cmd_ready        ;
  wire                arbt_bus_icb_cmd_sel          ;
  wire                arbt_bus_icb_cmd_read         ;
  wire    [  31:   0] arbt_bus_icb_cmd_addr         ;
  wire    [  63:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] arbt_bus_icb_cmd_size         ;
  wire                arbt_bus_icb_cmd_lock         ;
  wire                arbt_bus_icb_cmd_excl         ;
  wire    [   7:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] arbt_bus_icb_cmd_modes        ;
  wire                arbt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] arbt_bus_icb_cmd_attri        ;
  wire    [   1:   0] arbt_bus_icb_cmd_beat         ;
  wire    [   2:   0] arbt_bus_icb_cmd_usr          ;
  wire                arbt_bus_icb_rsp_ready        ;
  wire                arbt_bus_icb_rsp_valid        ;
  wire                arbt_bus_icb_rsp_err          ;
  wire                arbt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i0_icb_cmd_usr
                           };
      assign                 { i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (1),
  .ARBT_PTR_W (1),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid                   ),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready                   ),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read                    ),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [  31:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [  63:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [   7:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [   2:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock                    ),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl                    ),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [   7:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [   1:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [   1:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode                   ),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [   2:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [   1:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [   2:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready                   ),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid                   ),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err                     ),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok                 ),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [  63:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [   2:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_mgrp6_ficbnto1_bus #(
  parameter SUPPORT_LOCK = 1,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter ARBT_FIFO_OUTS_NUM    = 1,
  parameter ARBT_FIFO_OUTS_CNT_W  = 1,
  parameter ARBT_FIFO_CUT_READY   = 1,
  parameter RRBIN_CUT_TIMING = 0,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_ALLOW_0CYCL_RSP = 0
)(
  output icbnto1_active,
  input  i_clk_en,
  input  o_clk_en,
    output             o_icb_cmd_valid               ,
  input              o_icb_cmd_ready               ,
  output             o_icb_cmd_sel                 ,
  output             o_icb_cmd_read                ,
  output [  31:   0] o_icb_cmd_addr                ,
  output [  63:   0] o_icb_cmd_wdata               ,
  output [   7:   0] o_icb_cmd_wmask               ,
  output [   2:   0] o_icb_cmd_size                ,
  output             o_icb_cmd_lock                ,
  output             o_icb_cmd_excl                ,
  output [   7:   0] o_icb_cmd_xlen                ,
  output [   1:   0] o_icb_cmd_xburst              ,
  output [   1:   0] o_icb_cmd_modes               ,
  output             o_icb_cmd_dmode               ,
  output [   2:   0] o_icb_cmd_attri               ,
  output [   1:   0] o_icb_cmd_beat                ,
  output [   2:   0] o_icb_cmd_usr                 ,
  output             o_icb_rsp_ready               ,
  input              o_icb_rsp_valid               ,
  input              o_icb_rsp_err                 ,
  input              o_icb_rsp_excl_ok             ,
  input  [  63:   0] o_icb_rsp_rdata               ,
  input  [   2:   0] o_icb_rsp_usr                 ,
    input              i0_icb_cmd_valid              ,
  output             i0_icb_cmd_ready              ,
  input              i0_icb_cmd_sel                ,
  input              i0_icb_cmd_read               ,
  input  [  31:   0] i0_icb_cmd_addr               ,
  input  [  63:   0] i0_icb_cmd_wdata              ,
  input  [   7:   0] i0_icb_cmd_wmask              ,
  input  [   2:   0] i0_icb_cmd_size               ,
  input              i0_icb_cmd_lock               ,
  input              i0_icb_cmd_excl               ,
  input  [   7:   0] i0_icb_cmd_xlen               ,
  input  [   1:   0] i0_icb_cmd_xburst             ,
  input  [   1:   0] i0_icb_cmd_modes              ,
  input              i0_icb_cmd_dmode              ,
  input  [   2:   0] i0_icb_cmd_attri              ,
  input  [   1:   0] i0_icb_cmd_beat               ,
  input  [   2:   0] i0_icb_cmd_usr                ,
  input              i0_icb_rsp_ready              ,
  output             i0_icb_rsp_valid              ,
  output             i0_icb_rsp_err                ,
  output             i0_icb_rsp_excl_ok            ,
  output [  63:   0] i0_icb_rsp_rdata              ,
  output [   2:   0] i0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                arbt_bus_icb_cmd_valid        ;
  wire                arbt_bus_icb_cmd_ready        ;
  wire                arbt_bus_icb_cmd_sel          ;
  wire                arbt_bus_icb_cmd_read         ;
  wire    [  31:   0] arbt_bus_icb_cmd_addr         ;
  wire    [  63:   0] arbt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] arbt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] arbt_bus_icb_cmd_size         ;
  wire                arbt_bus_icb_cmd_lock         ;
  wire                arbt_bus_icb_cmd_excl         ;
  wire    [   7:   0] arbt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] arbt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] arbt_bus_icb_cmd_modes        ;
  wire                arbt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] arbt_bus_icb_cmd_attri        ;
  wire    [   1:   0] arbt_bus_icb_cmd_beat         ;
  wire    [   2:   0] arbt_bus_icb_cmd_usr          ;
  wire                arbt_bus_icb_rsp_ready        ;
  wire                arbt_bus_icb_rsp_valid        ;
  wire                arbt_bus_icb_rsp_err          ;
  wire                arbt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] arbt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] arbt_bus_icb_rsp_usr          ;
    assign arbt_bus_icb_cmd_valid =
                           { i0_icb_cmd_valid
                           };
    assign arbt_bus_icb_cmd_sel =
                           { i0_icb_cmd_sel
                           };
    assign arbt_bus_icb_cmd_read =
                           { i0_icb_cmd_read
                           };
    assign arbt_bus_icb_cmd_addr =
                           { i0_icb_cmd_addr
                           };
    assign arbt_bus_icb_cmd_wdata =
                           { i0_icb_cmd_wdata
                           };
    assign arbt_bus_icb_cmd_wmask =
                           { i0_icb_cmd_wmask
                           };
    assign arbt_bus_icb_cmd_size =
                           { i0_icb_cmd_size
                           };
    assign arbt_bus_icb_cmd_lock =
                           { i0_icb_cmd_lock
                           };
    assign arbt_bus_icb_cmd_excl =
                           { i0_icb_cmd_excl
                           };
    assign arbt_bus_icb_cmd_xlen =
                           { i0_icb_cmd_xlen
                           };
    assign arbt_bus_icb_cmd_xburst =
                           { i0_icb_cmd_xburst
                           };
    assign arbt_bus_icb_cmd_modes =
                           { i0_icb_cmd_modes
                           };
    assign arbt_bus_icb_cmd_dmode =
                           { i0_icb_cmd_dmode
                           };
    assign arbt_bus_icb_cmd_attri =
                           { i0_icb_cmd_attri
                           };
    assign arbt_bus_icb_cmd_beat =
                           { i0_icb_cmd_beat
                           };
    assign arbt_bus_icb_cmd_usr =
                           { i0_icb_cmd_usr
                           };
      assign                 { i0_icb_cmd_ready
                           } = arbt_bus_icb_cmd_ready;
      assign                 { i0_icb_rsp_valid
                           } = arbt_bus_icb_rsp_valid;
      assign                 { i0_icb_rsp_err
                           } = arbt_bus_icb_rsp_err;
      assign                 { i0_icb_rsp_excl_ok
                           } = arbt_bus_icb_rsp_excl_ok;
      assign                 { i0_icb_rsp_rdata
                           } = arbt_bus_icb_rsp_rdata;
      assign                 { i0_icb_rsp_usr
                           } = arbt_bus_icb_rsp_usr;
    assign arbt_bus_icb_rsp_ready =
                           { i0_icb_rsp_ready
                           };
    wire                arbt_icb_cmd_valid            ;
  wire                arbt_icb_cmd_ready            ;
  wire                arbt_icb_cmd_sel              ;
  wire                arbt_icb_cmd_read             ;
  wire    [  31:   0] arbt_icb_cmd_addr             ;
  wire    [  63:   0] arbt_icb_cmd_wdata            ;
  wire    [   7:   0] arbt_icb_cmd_wmask            ;
  wire    [   2:   0] arbt_icb_cmd_size             ;
  wire                arbt_icb_cmd_lock             ;
  wire                arbt_icb_cmd_excl             ;
  wire    [   7:   0] arbt_icb_cmd_xlen             ;
  wire    [   1:   0] arbt_icb_cmd_xburst           ;
  wire    [   1:   0] arbt_icb_cmd_modes            ;
  wire                arbt_icb_cmd_dmode            ;
  wire    [   2:   0] arbt_icb_cmd_attri            ;
  wire    [   1:   0] arbt_icb_cmd_beat             ;
  wire    [   2:   0] arbt_icb_cmd_usr              ;
  wire                arbt_icb_rsp_ready            ;
  wire                arbt_icb_rsp_valid            ;
  wire                arbt_icb_rsp_err              ;
  wire                arbt_icb_rsp_excl_ok          ;
  wire    [  63:   0] arbt_icb_rsp_rdata            ;
  wire    [   2:   0] arbt_icb_rsp_usr              ;
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire arbt_active;
  e603_subsys_gnrl_ficb_arbt # (
  .SUPPORT_LOCK(SUPPORT_LOCK),
  .ARBT_SCHEME (ARBT_SCHEME),
  .RRBIN_CUT_TIMING(RRBIN_CUT_TIMING),
    .PAYLOAD_NORST(PAYLOAD_NORST),
  .ALLOW_0CYCL_RSP (ARBT_ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (ARBT_FIFO_OUTS_NUM),
  .FIFO_CUT_READY  (ARBT_FIFO_CUT_READY),
  .ARBT_NUM   (1),
  .ARBT_PTR_W (1),
  .CMD_UW      (3),
  .RSP_UW      (3),
  .AW         (32),
  .DW         (64) 
  ) u_icb_arbt(
  .clk_en(i_clk_en),
  .arbt_active            (arbt_active),
      .i_bus_icb_cmd_valid            (arbt_bus_icb_cmd_valid                   ),
  .i_bus_icb_cmd_ready            (arbt_bus_icb_cmd_ready                   ),
  .i_bus_icb_cmd_read             (arbt_bus_icb_cmd_read                    ),
  .i_bus_icb_cmd_addr             (arbt_bus_icb_cmd_addr         [  31:   0]),
  .i_bus_icb_cmd_wdata            (arbt_bus_icb_cmd_wdata        [  63:   0]),
  .i_bus_icb_cmd_wmask            (arbt_bus_icb_cmd_wmask        [   7:   0]),
  .i_bus_icb_cmd_size             (arbt_bus_icb_cmd_size         [   2:   0]),
  .i_bus_icb_cmd_lock             (arbt_bus_icb_cmd_lock                    ),
  .i_bus_icb_cmd_excl             (arbt_bus_icb_cmd_excl                    ),
  .i_bus_icb_cmd_xlen             (arbt_bus_icb_cmd_xlen         [   7:   0]),
  .i_bus_icb_cmd_xburst           (arbt_bus_icb_cmd_xburst       [   1:   0]),
  .i_bus_icb_cmd_modes            (arbt_bus_icb_cmd_modes        [   1:   0]),
  .i_bus_icb_cmd_dmode            (arbt_bus_icb_cmd_dmode                   ),
  .i_bus_icb_cmd_attri            (arbt_bus_icb_cmd_attri        [   2:   0]),
  .i_bus_icb_cmd_beat             (arbt_bus_icb_cmd_beat         [   1:   0]),
  .i_bus_icb_cmd_usr              (arbt_bus_icb_cmd_usr          [   2:   0]),
  .i_bus_icb_rsp_ready            (arbt_bus_icb_rsp_ready                   ),
  .i_bus_icb_rsp_valid            (arbt_bus_icb_rsp_valid                   ),
  .i_bus_icb_rsp_err              (arbt_bus_icb_rsp_err                     ),
  .i_bus_icb_rsp_excl_ok          (arbt_bus_icb_rsp_excl_ok                 ),
  .i_bus_icb_rsp_rdata            (arbt_bus_icb_rsp_rdata        [  63:   0]),
  .i_bus_icb_rsp_usr              (arbt_bus_icb_rsp_usr          [   2:   0]),
      .o_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .o_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .o_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .o_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .o_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .o_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .o_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .o_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .o_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .o_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .o_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .o_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .o_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .o_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .o_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .o_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .o_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .o_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .o_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .o_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .o_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .o_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .o_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
    .i_bus_icb_cmd_sel_vec      (arbt_bus_icb_cmd_sel ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  wire buffer_active;
  assign icbnto1_active = buffer_active | arbt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (ARBT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (arbt_icb_cmd_valid                       ),
  .i_icb_cmd_ready                (arbt_icb_cmd_ready                       ),
  .i_icb_cmd_sel                  (arbt_icb_cmd_sel                         ),
  .i_icb_cmd_read                 (arbt_icb_cmd_read                        ),
  .i_icb_cmd_addr                 (arbt_icb_cmd_addr             [  31:   0]),
  .i_icb_cmd_wdata                (arbt_icb_cmd_wdata            [  63:   0]),
  .i_icb_cmd_wmask                (arbt_icb_cmd_wmask            [   7:   0]),
  .i_icb_cmd_size                 (arbt_icb_cmd_size             [   2:   0]),
  .i_icb_cmd_lock                 (arbt_icb_cmd_lock                        ),
  .i_icb_cmd_excl                 (arbt_icb_cmd_excl                        ),
  .i_icb_cmd_xlen                 (arbt_icb_cmd_xlen             [   7:   0]),
  .i_icb_cmd_xburst               (arbt_icb_cmd_xburst           [   1:   0]),
  .i_icb_cmd_modes                (arbt_icb_cmd_modes            [   1:   0]),
  .i_icb_cmd_dmode                (arbt_icb_cmd_dmode                       ),
  .i_icb_cmd_attri                (arbt_icb_cmd_attri            [   2:   0]),
  .i_icb_cmd_beat                 (arbt_icb_cmd_beat             [   1:   0]),
  .i_icb_cmd_usr                  (arbt_icb_cmd_usr              [   2:   0]),
  .i_icb_rsp_ready                (arbt_icb_rsp_ready                       ),
  .i_icb_rsp_valid                (arbt_icb_rsp_valid                       ),
  .i_icb_rsp_err                  (arbt_icb_rsp_err                         ),
  .i_icb_rsp_excl_ok              (arbt_icb_rsp_excl_ok                     ),
  .i_icb_rsp_rdata                (arbt_icb_rsp_rdata            [  63:   0]),
  .i_icb_rsp_usr                  (arbt_icb_rsp_usr              [   2:   0]),
      .o_icb_cmd_valid                (o_icb_cmd_valid                          ),
  .o_icb_cmd_ready                (o_icb_cmd_ready                          ),
  .o_icb_cmd_sel                  (o_icb_cmd_sel                            ),
  .o_icb_cmd_read                 (o_icb_cmd_read                           ),
  .o_icb_cmd_addr                 (o_icb_cmd_addr                [  31:   0]),
  .o_icb_cmd_wdata                (o_icb_cmd_wdata               [  63:   0]),
  .o_icb_cmd_wmask                (o_icb_cmd_wmask               [   7:   0]),
  .o_icb_cmd_size                 (o_icb_cmd_size                [   2:   0]),
  .o_icb_cmd_lock                 (o_icb_cmd_lock                           ),
  .o_icb_cmd_excl                 (o_icb_cmd_excl                           ),
  .o_icb_cmd_xlen                 (o_icb_cmd_xlen                [   7:   0]),
  .o_icb_cmd_xburst               (o_icb_cmd_xburst              [   1:   0]),
  .o_icb_cmd_modes                (o_icb_cmd_modes               [   1:   0]),
  .o_icb_cmd_dmode                (o_icb_cmd_dmode                          ),
  .o_icb_cmd_attri                (o_icb_cmd_attri               [   2:   0]),
  .o_icb_cmd_beat                 (o_icb_cmd_beat                [   1:   0]),
  .o_icb_cmd_usr                  (o_icb_cmd_usr                 [   2:   0]),
  .o_icb_rsp_ready                (o_icb_rsp_ready                          ),
  .o_icb_rsp_valid                (o_icb_rsp_valid                          ),
  .o_icb_rsp_err                  (o_icb_rsp_err                            ),
  .o_icb_rsp_excl_ok              (o_icb_rsp_excl_ok                        ),
  .o_icb_rsp_rdata                (o_icb_rsp_rdata               [  63:   0]),
  .o_icb_rsp_usr                  (o_icb_rsp_usr                 [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
endmodule
module e603_subsys_sgrp0_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
        wire                o1_icb_cmd_valid              ;
  wire                o1_icb_cmd_ready              ;
  wire                o1_icb_cmd_sel                ;
  wire                o1_icb_cmd_read               ;
  wire    [  31:   0] o1_icb_cmd_addr               ;
  wire    [  63:   0] o1_icb_cmd_wdata              ;
  wire    [   7:   0] o1_icb_cmd_wmask              ;
  wire    [   2:   0] o1_icb_cmd_size               ;
  wire                o1_icb_cmd_lock               ;
  wire                o1_icb_cmd_excl               ;
  wire    [   7:   0] o1_icb_cmd_xlen               ;
  wire    [   1:   0] o1_icb_cmd_xburst             ;
  wire    [   1:   0] o1_icb_cmd_modes              ;
  wire                o1_icb_cmd_dmode              ;
  wire    [   2:   0] o1_icb_cmd_attri              ;
  wire    [   1:   0] o1_icb_cmd_beat               ;
  wire    [   2:   0] o1_icb_cmd_usr                ;
  wire                o1_icb_rsp_ready              ;
  wire                o1_icb_rsp_valid              ;
  wire                o1_icb_rsp_err                ;
  wire                o1_icb_rsp_excl_ok            ;
  wire    [  63:   0] o1_icb_rsp_rdata              ;
  wire    [   2:   0] o1_icb_rsp_usr                ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_read                 (i_icb_cmd_read                           ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   1:   0] splt_bus_icb_cmd_valid        ;
  wire    [   1:   0] splt_bus_icb_cmd_ready        ;
  wire    [   1:   0] splt_bus_icb_cmd_sel          ;
  wire    [   1:   0] splt_bus_icb_cmd_read         ;
  wire    [  63:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 127:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  15:   0] splt_bus_icb_cmd_wmask        ;
  wire    [   5:   0] splt_bus_icb_cmd_size         ;
  wire    [   1:   0] splt_bus_icb_cmd_lock         ;
  wire    [   1:   0] splt_bus_icb_cmd_excl         ;
  wire    [  15:   0] splt_bus_icb_cmd_xlen         ;
  wire    [   3:   0] splt_bus_icb_cmd_xburst       ;
  wire    [   3:   0] splt_bus_icb_cmd_modes        ;
  wire    [   1:   0] splt_bus_icb_cmd_dmode        ;
  wire    [   5:   0] splt_bus_icb_cmd_attri        ;
  wire    [   3:   0] splt_bus_icb_cmd_beat         ;
  wire    [   5:   0] splt_bus_icb_cmd_usr          ;
  wire    [   1:   0] splt_bus_icb_rsp_ready        ;
  wire    [   1:   0] splt_bus_icb_rsp_valid        ;
  wire    [   1:   0] splt_bus_icb_rsp_err          ;
  wire    [   1:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 127:   0] splt_bus_icb_rsp_rdata        ;
  wire    [   5:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = 1'b1
                          & (~icb_cmd_o0)
                        ; 
  wire [2-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (2),
  .SPLT_PTR_W (2),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   1:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   1:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   1:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   1:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [  63:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 127:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  15:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [   5:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   1:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   1:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  15:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [   3:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [   3:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   1:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [   5:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [   3:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [   5:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   1:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   1:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   1:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   1:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 127:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [   5:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  assign  o1_icb_rsp_err     = 1'b1;
  assign  o1_icb_rsp_excl_ok = 1'b0;
  assign  o1_icb_rsp_rdata   = {64{1'b0}};
  assign  o1_icb_rsp_usr     = {3{1'b0}};
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_dft_rsp_gen_stage(
    .i_vld(o1_icb_cmd_valid & o_clk_en), 
    .i_rdy(o1_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(o1_icb_rsp_valid), 
    .o_rdy(o1_icb_rsp_ready & o_clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_sgrp1_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
        wire                o1_icb_cmd_valid              ;
  wire                o1_icb_cmd_ready              ;
  wire                o1_icb_cmd_sel                ;
  wire                o1_icb_cmd_read               ;
  wire    [  31:   0] o1_icb_cmd_addr               ;
  wire    [  63:   0] o1_icb_cmd_wdata              ;
  wire    [   7:   0] o1_icb_cmd_wmask              ;
  wire    [   2:   0] o1_icb_cmd_size               ;
  wire                o1_icb_cmd_lock               ;
  wire                o1_icb_cmd_excl               ;
  wire    [   7:   0] o1_icb_cmd_xlen               ;
  wire    [   1:   0] o1_icb_cmd_xburst             ;
  wire    [   1:   0] o1_icb_cmd_modes              ;
  wire                o1_icb_cmd_dmode              ;
  wire    [   2:   0] o1_icb_cmd_attri              ;
  wire    [   1:   0] o1_icb_cmd_beat               ;
  wire    [   2:   0] o1_icb_cmd_usr                ;
  wire                o1_icb_rsp_ready              ;
  wire                o1_icb_rsp_valid              ;
  wire                o1_icb_rsp_err                ;
  wire                o1_icb_rsp_excl_ok            ;
  wire    [  63:   0] o1_icb_rsp_rdata              ;
  wire    [   2:   0] o1_icb_rsp_usr                ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_read                 (i_icb_cmd_read                           ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   1:   0] splt_bus_icb_cmd_valid        ;
  wire    [   1:   0] splt_bus_icb_cmd_ready        ;
  wire    [   1:   0] splt_bus_icb_cmd_sel          ;
  wire    [   1:   0] splt_bus_icb_cmd_read         ;
  wire    [  63:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 127:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  15:   0] splt_bus_icb_cmd_wmask        ;
  wire    [   5:   0] splt_bus_icb_cmd_size         ;
  wire    [   1:   0] splt_bus_icb_cmd_lock         ;
  wire    [   1:   0] splt_bus_icb_cmd_excl         ;
  wire    [  15:   0] splt_bus_icb_cmd_xlen         ;
  wire    [   3:   0] splt_bus_icb_cmd_xburst       ;
  wire    [   3:   0] splt_bus_icb_cmd_modes        ;
  wire    [   1:   0] splt_bus_icb_cmd_dmode        ;
  wire    [   5:   0] splt_bus_icb_cmd_attri        ;
  wire    [   3:   0] splt_bus_icb_cmd_beat         ;
  wire    [   5:   0] splt_bus_icb_cmd_usr          ;
  wire    [   1:   0] splt_bus_icb_rsp_ready        ;
  wire    [   1:   0] splt_bus_icb_rsp_valid        ;
  wire    [   1:   0] splt_bus_icb_rsp_err          ;
  wire    [   1:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 127:   0] splt_bus_icb_rsp_rdata        ;
  wire    [   5:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = 1'b1
                          & (~icb_cmd_o0)
                        ; 
  wire [2-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (2),
  .SPLT_PTR_W (2),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   1:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   1:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   1:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   1:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [  63:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 127:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  15:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [   5:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   1:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   1:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  15:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [   3:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [   3:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   1:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [   5:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [   3:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [   5:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   1:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   1:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   1:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   1:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 127:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [   5:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  assign  o1_icb_rsp_err     = 1'b1;
  assign  o1_icb_rsp_excl_ok = 1'b0;
  assign  o1_icb_rsp_rdata   = {64{1'b0}};
  assign  o1_icb_rsp_usr     = {3{1'b0}};
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_dft_rsp_gen_stage(
    .i_vld(o1_icb_cmd_valid & o_clk_en), 
    .i_rdy(o1_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(o1_icb_rsp_valid), 
    .o_rdy(o1_icb_rsp_ready & o_clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_sgrp2_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
        wire                o1_icb_cmd_valid              ;
  wire                o1_icb_cmd_ready              ;
  wire                o1_icb_cmd_sel                ;
  wire                o1_icb_cmd_read               ;
  wire    [  31:   0] o1_icb_cmd_addr               ;
  wire    [  63:   0] o1_icb_cmd_wdata              ;
  wire    [   7:   0] o1_icb_cmd_wmask              ;
  wire    [   2:   0] o1_icb_cmd_size               ;
  wire                o1_icb_cmd_lock               ;
  wire                o1_icb_cmd_excl               ;
  wire    [   7:   0] o1_icb_cmd_xlen               ;
  wire    [   1:   0] o1_icb_cmd_xburst             ;
  wire    [   1:   0] o1_icb_cmd_modes              ;
  wire                o1_icb_cmd_dmode              ;
  wire    [   2:   0] o1_icb_cmd_attri              ;
  wire    [   1:   0] o1_icb_cmd_beat               ;
  wire    [   2:   0] o1_icb_cmd_usr                ;
  wire                o1_icb_rsp_ready              ;
  wire                o1_icb_rsp_valid              ;
  wire                o1_icb_rsp_err                ;
  wire                o1_icb_rsp_excl_ok            ;
  wire    [  63:   0] o1_icb_rsp_rdata              ;
  wire    [   2:   0] o1_icb_rsp_usr                ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_read                 (i_icb_cmd_read                           ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   1:   0] splt_bus_icb_cmd_valid        ;
  wire    [   1:   0] splt_bus_icb_cmd_ready        ;
  wire    [   1:   0] splt_bus_icb_cmd_sel          ;
  wire    [   1:   0] splt_bus_icb_cmd_read         ;
  wire    [  63:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 127:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  15:   0] splt_bus_icb_cmd_wmask        ;
  wire    [   5:   0] splt_bus_icb_cmd_size         ;
  wire    [   1:   0] splt_bus_icb_cmd_lock         ;
  wire    [   1:   0] splt_bus_icb_cmd_excl         ;
  wire    [  15:   0] splt_bus_icb_cmd_xlen         ;
  wire    [   3:   0] splt_bus_icb_cmd_xburst       ;
  wire    [   3:   0] splt_bus_icb_cmd_modes        ;
  wire    [   1:   0] splt_bus_icb_cmd_dmode        ;
  wire    [   5:   0] splt_bus_icb_cmd_attri        ;
  wire    [   3:   0] splt_bus_icb_cmd_beat         ;
  wire    [   5:   0] splt_bus_icb_cmd_usr          ;
  wire    [   1:   0] splt_bus_icb_rsp_ready        ;
  wire    [   1:   0] splt_bus_icb_rsp_valid        ;
  wire    [   1:   0] splt_bus_icb_rsp_err          ;
  wire    [   1:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 127:   0] splt_bus_icb_rsp_rdata        ;
  wire    [   5:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = 1'b1
                          & (~icb_cmd_o0)
                        ; 
  wire [2-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (2),
  .SPLT_PTR_W (2),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   1:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   1:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   1:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   1:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [  63:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 127:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  15:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [   5:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   1:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   1:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  15:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [   3:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [   3:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   1:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [   5:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [   3:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [   5:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   1:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   1:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   1:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   1:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 127:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [   5:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  assign  o1_icb_rsp_err     = 1'b1;
  assign  o1_icb_rsp_excl_ok = 1'b0;
  assign  o1_icb_rsp_rdata   = {64{1'b0}};
  assign  o1_icb_rsp_usr     = {3{1'b0}};
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_dft_rsp_gen_stage(
    .i_vld(o1_icb_cmd_valid & o_clk_en), 
    .i_rdy(o1_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(o1_icb_rsp_valid), 
    .o_rdy(o1_icb_rsp_ready & o_clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_sgrp3_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
        wire                o1_icb_cmd_valid              ;
  wire                o1_icb_cmd_ready              ;
  wire                o1_icb_cmd_sel                ;
  wire                o1_icb_cmd_read               ;
  wire    [  31:   0] o1_icb_cmd_addr               ;
  wire    [  63:   0] o1_icb_cmd_wdata              ;
  wire    [   7:   0] o1_icb_cmd_wmask              ;
  wire    [   2:   0] o1_icb_cmd_size               ;
  wire                o1_icb_cmd_lock               ;
  wire                o1_icb_cmd_excl               ;
  wire    [   7:   0] o1_icb_cmd_xlen               ;
  wire    [   1:   0] o1_icb_cmd_xburst             ;
  wire    [   1:   0] o1_icb_cmd_modes              ;
  wire                o1_icb_cmd_dmode              ;
  wire    [   2:   0] o1_icb_cmd_attri              ;
  wire    [   1:   0] o1_icb_cmd_beat               ;
  wire    [   2:   0] o1_icb_cmd_usr                ;
  wire                o1_icb_rsp_ready              ;
  wire                o1_icb_rsp_valid              ;
  wire                o1_icb_rsp_err                ;
  wire                o1_icb_rsp_excl_ok            ;
  wire    [  63:   0] o1_icb_rsp_rdata              ;
  wire    [   2:   0] o1_icb_rsp_usr                ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_read                 (i_icb_cmd_read                           ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   1:   0] splt_bus_icb_cmd_valid        ;
  wire    [   1:   0] splt_bus_icb_cmd_ready        ;
  wire    [   1:   0] splt_bus_icb_cmd_sel          ;
  wire    [   1:   0] splt_bus_icb_cmd_read         ;
  wire    [  63:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 127:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  15:   0] splt_bus_icb_cmd_wmask        ;
  wire    [   5:   0] splt_bus_icb_cmd_size         ;
  wire    [   1:   0] splt_bus_icb_cmd_lock         ;
  wire    [   1:   0] splt_bus_icb_cmd_excl         ;
  wire    [  15:   0] splt_bus_icb_cmd_xlen         ;
  wire    [   3:   0] splt_bus_icb_cmd_xburst       ;
  wire    [   3:   0] splt_bus_icb_cmd_modes        ;
  wire    [   1:   0] splt_bus_icb_cmd_dmode        ;
  wire    [   5:   0] splt_bus_icb_cmd_attri        ;
  wire    [   3:   0] splt_bus_icb_cmd_beat         ;
  wire    [   5:   0] splt_bus_icb_cmd_usr          ;
  wire    [   1:   0] splt_bus_icb_rsp_ready        ;
  wire    [   1:   0] splt_bus_icb_rsp_valid        ;
  wire    [   1:   0] splt_bus_icb_rsp_err          ;
  wire    [   1:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 127:   0] splt_bus_icb_rsp_rdata        ;
  wire    [   5:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = 1'b1
                          & (~icb_cmd_o0)
                        ; 
  wire [2-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (2),
  .SPLT_PTR_W (2),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   1:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   1:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   1:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   1:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [  63:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 127:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  15:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [   5:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   1:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   1:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  15:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [   3:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [   3:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   1:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [   5:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [   3:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [   5:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   1:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   1:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   1:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   1:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 127:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [   5:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  assign  o1_icb_rsp_err     = 1'b1;
  assign  o1_icb_rsp_excl_ok = 1'b0;
  assign  o1_icb_rsp_rdata   = {64{1'b0}};
  assign  o1_icb_rsp_usr     = {3{1'b0}};
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_dft_rsp_gen_stage(
    .i_vld(o1_icb_cmd_valid & o_clk_en), 
    .i_rdy(o1_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(o1_icb_rsp_valid), 
    .o_rdy(o1_icb_rsp_ready & o_clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_sgrp4_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter O2_BASE_ADDR       = 32'h0,       
  parameter O2_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input                          o1_icb_enable,
    output             o1_icb_cmd_valid              ,
  input              o1_icb_cmd_ready              ,
  output             o1_icb_cmd_sel                ,
  output             o1_icb_cmd_read               ,
  output [  31:   0] o1_icb_cmd_addr               ,
  output [  63:   0] o1_icb_cmd_wdata              ,
  output [   7:   0] o1_icb_cmd_wmask              ,
  output [   2:   0] o1_icb_cmd_size               ,
  output             o1_icb_cmd_lock               ,
  output             o1_icb_cmd_excl               ,
  output [   7:   0] o1_icb_cmd_xlen               ,
  output [   1:   0] o1_icb_cmd_xburst             ,
  output [   1:   0] o1_icb_cmd_modes              ,
  output             o1_icb_cmd_dmode              ,
  output [   2:   0] o1_icb_cmd_attri              ,
  output [   1:   0] o1_icb_cmd_beat               ,
  output [   2:   0] o1_icb_cmd_usr                ,
  output             o1_icb_rsp_ready              ,
  input              o1_icb_rsp_valid              ,
  input              o1_icb_rsp_err                ,
  input              o1_icb_rsp_excl_ok            ,
  input  [  63:   0] o1_icb_rsp_rdata              ,
  input  [   2:   0] o1_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
        wire                o2_icb_cmd_valid              ;
  wire                o2_icb_cmd_ready              ;
  wire                o2_icb_cmd_sel                ;
  wire                o2_icb_cmd_read               ;
  wire    [  31:   0] o2_icb_cmd_addr               ;
  wire    [  63:   0] o2_icb_cmd_wdata              ;
  wire    [   7:   0] o2_icb_cmd_wmask              ;
  wire    [   2:   0] o2_icb_cmd_size               ;
  wire                o2_icb_cmd_lock               ;
  wire                o2_icb_cmd_excl               ;
  wire    [   7:   0] o2_icb_cmd_xlen               ;
  wire    [   1:   0] o2_icb_cmd_xburst             ;
  wire    [   1:   0] o2_icb_cmd_modes              ;
  wire                o2_icb_cmd_dmode              ;
  wire    [   2:   0] o2_icb_cmd_attri              ;
  wire    [   1:   0] o2_icb_cmd_beat               ;
  wire    [   2:   0] o2_icb_cmd_usr                ;
  wire                o2_icb_rsp_ready              ;
  wire                o2_icb_rsp_valid              ;
  wire                o2_icb_rsp_err                ;
  wire                o2_icb_rsp_excl_ok            ;
  wire    [  63:   0] o2_icb_rsp_rdata              ;
  wire    [   2:   0] o2_icb_rsp_usr                ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_read                 (i_icb_cmd_read                           ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   2:   0] splt_bus_icb_cmd_valid        ;
  wire    [   2:   0] splt_bus_icb_cmd_ready        ;
  wire    [   2:   0] splt_bus_icb_cmd_sel          ;
  wire    [   2:   0] splt_bus_icb_cmd_read         ;
  wire    [  95:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 191:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  23:   0] splt_bus_icb_cmd_wmask        ;
  wire    [   8:   0] splt_bus_icb_cmd_size         ;
  wire    [   2:   0] splt_bus_icb_cmd_lock         ;
  wire    [   2:   0] splt_bus_icb_cmd_excl         ;
  wire    [  23:   0] splt_bus_icb_cmd_xlen         ;
  wire    [   5:   0] splt_bus_icb_cmd_xburst       ;
  wire    [   5:   0] splt_bus_icb_cmd_modes        ;
  wire    [   2:   0] splt_bus_icb_cmd_dmode        ;
  wire    [   8:   0] splt_bus_icb_cmd_attri        ;
  wire    [   5:   0] splt_bus_icb_cmd_beat         ;
  wire    [   8:   0] splt_bus_icb_cmd_usr          ;
  wire    [   2:   0] splt_bus_icb_rsp_ready        ;
  wire    [   2:   0] splt_bus_icb_rsp_valid        ;
  wire    [   2:   0] splt_bus_icb_rsp_err          ;
  wire    [   2:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 191:   0] splt_bus_icb_rsp_rdata        ;
  wire    [   8:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o2_icb_cmd_sel
                           , o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o2_icb_cmd_valid
                           , o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o2_icb_cmd_read
                           , o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o2_icb_cmd_addr
                           , o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o2_icb_cmd_wdata
                           , o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o2_icb_cmd_wmask
                           , o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o2_icb_cmd_size
                           , o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o2_icb_cmd_lock
                           , o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o2_icb_cmd_excl
                           , o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o2_icb_cmd_xlen
                           , o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o2_icb_cmd_xburst
                           , o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o2_icb_cmd_modes
                           , o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o2_icb_cmd_dmode
                           , o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o2_icb_cmd_attri
                           , o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o2_icb_cmd_beat
                           , o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o2_icb_cmd_usr
                           , o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o2_icb_cmd_ready
                           , o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o2_icb_rsp_valid
                           , o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o2_icb_rsp_err
                           , o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o2_icb_rsp_excl_ok
                           , o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o2_icb_rsp_rdata
                           , o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o2_icb_rsp_usr
                           , o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o2_icb_rsp_ready
                           , o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = (buf_icb_cmd_addr     [31:O1_BASE_REGION_LSB]
                         ==  O1_BASE_ADDR [31:O1_BASE_REGION_LSB] 
                        ) & o1_icb_enable 
                          & (~icb_cmd_o0)
                        ; 
      wire icb_cmd_o2 = 1'b1
                          & (~icb_cmd_o0)
                          & (~icb_cmd_o1)
                        ; 
  wire [3-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o2
                    , icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (3),
  .SPLT_PTR_W (3),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   2:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   2:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   2:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   2:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [  95:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 191:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  23:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [   8:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   2:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   2:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  23:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [   5:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [   5:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   2:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [   8:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [   5:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [   8:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   2:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   2:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   2:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   2:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 191:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [   8:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  assign  o2_icb_rsp_err     = 1'b1;
  assign  o2_icb_rsp_excl_ok = 1'b0;
  assign  o2_icb_rsp_rdata   = {64{1'b0}};
  assign  o2_icb_rsp_usr     = {3{1'b0}};
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_dft_rsp_gen_stage(
    .i_vld(o2_icb_cmd_valid & o_clk_en), 
    .i_rdy(o2_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(o2_icb_rsp_valid), 
    .o_rdy(o2_icb_rsp_ready & o_clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_sgrp5_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter O1_BASE_ADDR       = 32'h0,       
  parameter O1_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
  input                          o0_icb_enable,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
        wire                o1_icb_cmd_valid              ;
  wire                o1_icb_cmd_ready              ;
  wire                o1_icb_cmd_sel                ;
  wire                o1_icb_cmd_read               ;
  wire    [  31:   0] o1_icb_cmd_addr               ;
  wire    [  63:   0] o1_icb_cmd_wdata              ;
  wire    [   7:   0] o1_icb_cmd_wmask              ;
  wire    [   2:   0] o1_icb_cmd_size               ;
  wire                o1_icb_cmd_lock               ;
  wire                o1_icb_cmd_excl               ;
  wire    [   7:   0] o1_icb_cmd_xlen               ;
  wire    [   1:   0] o1_icb_cmd_xburst             ;
  wire    [   1:   0] o1_icb_cmd_modes              ;
  wire                o1_icb_cmd_dmode              ;
  wire    [   2:   0] o1_icb_cmd_attri              ;
  wire    [   1:   0] o1_icb_cmd_beat               ;
  wire    [   2:   0] o1_icb_cmd_usr                ;
  wire                o1_icb_rsp_ready              ;
  wire                o1_icb_rsp_valid              ;
  wire                o1_icb_rsp_err                ;
  wire                o1_icb_rsp_excl_ok            ;
  wire    [  63:   0] o1_icb_rsp_rdata              ;
  wire    [   2:   0] o1_icb_rsp_usr                ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(ICB_FIFO_CMD_BYPBUF),
    .CMD_DP(ICB_FIFO_CMD_DP),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_read                 (i_icb_cmd_read                           ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire    [   1:   0] splt_bus_icb_cmd_valid        ;
  wire    [   1:   0] splt_bus_icb_cmd_ready        ;
  wire    [   1:   0] splt_bus_icb_cmd_sel          ;
  wire    [   1:   0] splt_bus_icb_cmd_read         ;
  wire    [  63:   0] splt_bus_icb_cmd_addr         ;
  wire    [ 127:   0] splt_bus_icb_cmd_wdata        ;
  wire    [  15:   0] splt_bus_icb_cmd_wmask        ;
  wire    [   5:   0] splt_bus_icb_cmd_size         ;
  wire    [   1:   0] splt_bus_icb_cmd_lock         ;
  wire    [   1:   0] splt_bus_icb_cmd_excl         ;
  wire    [  15:   0] splt_bus_icb_cmd_xlen         ;
  wire    [   3:   0] splt_bus_icb_cmd_xburst       ;
  wire    [   3:   0] splt_bus_icb_cmd_modes        ;
  wire    [   1:   0] splt_bus_icb_cmd_dmode        ;
  wire    [   5:   0] splt_bus_icb_cmd_attri        ;
  wire    [   3:   0] splt_bus_icb_cmd_beat         ;
  wire    [   5:   0] splt_bus_icb_cmd_usr          ;
  wire    [   1:   0] splt_bus_icb_rsp_ready        ;
  wire    [   1:   0] splt_bus_icb_rsp_valid        ;
  wire    [   1:   0] splt_bus_icb_rsp_err          ;
  wire    [   1:   0] splt_bus_icb_rsp_excl_ok      ;
  wire    [ 127:   0] splt_bus_icb_rsp_rdata        ;
  wire    [   5:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o1_icb_cmd_sel
                           , o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o1_icb_cmd_valid
                           , o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o1_icb_cmd_read
                           , o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o1_icb_cmd_addr
                           , o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o1_icb_cmd_wdata
                           , o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o1_icb_cmd_wmask
                           , o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o1_icb_cmd_size
                           , o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o1_icb_cmd_lock
                           , o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o1_icb_cmd_excl
                           , o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o1_icb_cmd_xlen
                           , o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o1_icb_cmd_xburst
                           , o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o1_icb_cmd_modes
                           , o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o1_icb_cmd_dmode
                           , o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o1_icb_cmd_attri
                           , o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o1_icb_cmd_beat
                           , o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o1_icb_cmd_usr
                           , o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o1_icb_cmd_ready
                           , o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o1_icb_rsp_valid
                           , o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o1_icb_rsp_err
                           , o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o1_icb_rsp_excl_ok
                           , o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o1_icb_rsp_rdata
                           , o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o1_icb_rsp_usr
                           , o0_icb_rsp_usr
                           };
      assign                 { o1_icb_rsp_ready
                           , o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = (buf_icb_cmd_addr     [31:O0_BASE_REGION_LSB]
                         ==  O0_BASE_ADDR [31:O0_BASE_REGION_LSB] 
                        ) & o0_icb_enable 
                        ; 
      wire icb_cmd_o1 = 1'b1
                          & (~icb_cmd_o0)
                        ; 
  wire [2-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o1
                    , icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (2),
  .SPLT_PTR_W (2),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid        [   1:   0]),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready        [   1:   0]),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel          [   1:   0]),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read         [   1:   0]),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [  63:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [ 127:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [  15:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [   5:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock         [   1:   0]),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl         [   1:   0]),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [  15:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [   3:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [   3:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode        [   1:   0]),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [   5:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [   3:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [   5:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready        [   1:   0]),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid        [   1:   0]),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err          [   1:   0]),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok      [   1:   0]),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [ 127:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [   5:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
  assign  o1_icb_rsp_err     = 1'b1;
  assign  o1_icb_rsp_excl_ok = 1'b0;
  assign  o1_icb_rsp_rdata   = {64{1'b0}};
  assign  o1_icb_rsp_usr     = {3{1'b0}};
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_dft_rsp_gen_stage(
    .i_vld(o1_icb_cmd_valid & o_clk_en), 
    .i_rdy(o1_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(o1_icb_rsp_valid), 
    .o_rdy(o1_icb_rsp_ready & o_clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_sgrp6_ficb1ton_bus #(
  parameter I_SUPPORT_RATIO = 0, 
  parameter O_SUPPORT_RATIO = 0,
  parameter ALLOW_DIFF =0,
  parameter ALLOW_0CYCL_RSP =0,
  parameter ICB_FIFO_CMD_BYPBUF = 0,
  parameter ICB_FIFO_CMD_DP = 0, 
  parameter ICB_FIFO_RSP_DP = 0, 
  parameter ICB_FIFO_CMD_CUT_READY = 1, 
  parameter ICB_FIFO_RSP_CUT_READY = 1, 
  parameter O0_BASE_ADDR       = 32'h0,       
  parameter O0_BASE_REGION_LSB = 12,
  parameter PAYLOAD_NORST    = 0,
  parameter SPLT_FIFO_OUTS_NUM    = 1,
  parameter SPLT_FIFO_OUTS_CNT_W  = 1,
  parameter SPLT_FIFO_CUT_READY   = 1 
)(
  input i_clk_en,
  input o_clk_en,
  output  icb1ton_active,
    input              i_icb_cmd_valid               ,
  output             i_icb_cmd_ready               ,
  input              i_icb_cmd_sel                 ,
  input              i_icb_cmd_read                ,
  input  [  31:   0] i_icb_cmd_addr                ,
  input  [  63:   0] i_icb_cmd_wdata               ,
  input  [   7:   0] i_icb_cmd_wmask               ,
  input  [   2:   0] i_icb_cmd_size                ,
  input              i_icb_cmd_lock                ,
  input              i_icb_cmd_excl                ,
  input  [   7:   0] i_icb_cmd_xlen                ,
  input  [   1:   0] i_icb_cmd_xburst              ,
  input  [   1:   0] i_icb_cmd_modes               ,
  input              i_icb_cmd_dmode               ,
  input  [   2:   0] i_icb_cmd_attri               ,
  input  [   1:   0] i_icb_cmd_beat                ,
  input  [   2:   0] i_icb_cmd_usr                 ,
  input              i_icb_rsp_ready               ,
  output             i_icb_rsp_valid               ,
  output             i_icb_rsp_err                 ,
  output             i_icb_rsp_excl_ok             ,
  output [  63:   0] i_icb_rsp_rdata               ,
  output [   2:   0] i_icb_rsp_usr                 ,
    output             o0_icb_cmd_valid              ,
  input              o0_icb_cmd_ready              ,
  output             o0_icb_cmd_sel                ,
  output             o0_icb_cmd_read               ,
  output [  31:   0] o0_icb_cmd_addr               ,
  output [  63:   0] o0_icb_cmd_wdata              ,
  output [   7:   0] o0_icb_cmd_wmask              ,
  output [   2:   0] o0_icb_cmd_size               ,
  output             o0_icb_cmd_lock               ,
  output             o0_icb_cmd_excl               ,
  output [   7:   0] o0_icb_cmd_xlen               ,
  output [   1:   0] o0_icb_cmd_xburst             ,
  output [   1:   0] o0_icb_cmd_modes              ,
  output             o0_icb_cmd_dmode              ,
  output [   2:   0] o0_icb_cmd_attri              ,
  output [   1:   0] o0_icb_cmd_beat               ,
  output [   2:   0] o0_icb_cmd_usr                ,
  output             o0_icb_rsp_ready              ,
  input              o0_icb_rsp_valid              ,
  input              o0_icb_rsp_err                ,
  input              o0_icb_rsp_excl_ok            ,
  input  [  63:   0] o0_icb_rsp_rdata              ,
  input  [   2:   0] o0_icb_rsp_usr                ,
  input  clk,
  input  rst_n
  );
    wire                buf_icb_cmd_valid             ;
  wire                buf_icb_cmd_ready             ;
  wire                buf_icb_cmd_sel               ;
  wire                buf_icb_cmd_read              ;
  wire    [  31:   0] buf_icb_cmd_addr              ;
  wire    [  63:   0] buf_icb_cmd_wdata             ;
  wire    [   7:   0] buf_icb_cmd_wmask             ;
  wire    [   2:   0] buf_icb_cmd_size              ;
  wire                buf_icb_cmd_lock              ;
  wire                buf_icb_cmd_excl              ;
  wire    [   7:   0] buf_icb_cmd_xlen              ;
  wire    [   1:   0] buf_icb_cmd_xburst            ;
  wire    [   1:   0] buf_icb_cmd_modes             ;
  wire                buf_icb_cmd_dmode             ;
  wire    [   2:   0] buf_icb_cmd_attri             ;
  wire    [   1:   0] buf_icb_cmd_beat              ;
  wire    [   2:   0] buf_icb_cmd_usr               ;
  wire                buf_icb_rsp_ready             ;
  wire                buf_icb_rsp_valid             ;
  wire                buf_icb_rsp_err               ;
  wire                buf_icb_rsp_excl_ok           ;
  wire    [  63:   0] buf_icb_rsp_rdata             ;
  wire    [   2:   0] buf_icb_rsp_usr               ;
  wire buffer_active;
  wire splt_active;
  assign icb1ton_active = buffer_active | splt_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(I_SUPPORT_RATIO),
    .O_SUPPORT_RATIO(O_SUPPORT_RATIO),
    .OUTS_CNT_W     (SPLT_FIFO_OUTS_CNT_W),
    .AW    (32),
    .DW    (64), 
    .RSP_DP(ICB_FIFO_RSP_DP),
    .CMD_BYPBUF(0),
    .CMD_DP(0),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .CMD_CUT_READY (ICB_FIFO_CMD_CUT_READY),
    .RSP_CUT_READY (ICB_FIFO_RSP_CUT_READY),
    .CMD_UW (3),
    .RSP_UW (3)
  )u_e603_subsys_icb_buffer(
    .i_clk_en   (i_clk_en),
    .o_clk_en   (o_clk_en),
    .icb_buffer_active (buffer_active),
      .i_icb_cmd_valid                (i_icb_cmd_valid                          ),
  .i_icb_cmd_ready                (i_icb_cmd_ready                          ),
  .i_icb_cmd_sel                  (i_icb_cmd_sel                            ),
  .i_icb_cmd_read                 (i_icb_cmd_read                           ),
  .i_icb_cmd_addr                 (i_icb_cmd_addr                [  31:   0]),
  .i_icb_cmd_wdata                (i_icb_cmd_wdata               [  63:   0]),
  .i_icb_cmd_wmask                (i_icb_cmd_wmask               [   7:   0]),
  .i_icb_cmd_size                 (i_icb_cmd_size                [   2:   0]),
  .i_icb_cmd_lock                 (i_icb_cmd_lock                           ),
  .i_icb_cmd_excl                 (i_icb_cmd_excl                           ),
  .i_icb_cmd_xlen                 (i_icb_cmd_xlen                [   7:   0]),
  .i_icb_cmd_xburst               (i_icb_cmd_xburst              [   1:   0]),
  .i_icb_cmd_modes                (i_icb_cmd_modes               [   1:   0]),
  .i_icb_cmd_dmode                (i_icb_cmd_dmode                          ),
  .i_icb_cmd_attri                (i_icb_cmd_attri               [   2:   0]),
  .i_icb_cmd_beat                 (i_icb_cmd_beat                [   1:   0]),
  .i_icb_cmd_usr                  (i_icb_cmd_usr                 [   2:   0]),
  .i_icb_rsp_ready                (i_icb_rsp_ready                          ),
  .i_icb_rsp_valid                (i_icb_rsp_valid                          ),
  .i_icb_rsp_err                  (i_icb_rsp_err                            ),
  .i_icb_rsp_excl_ok              (i_icb_rsp_excl_ok                        ),
  .i_icb_rsp_rdata                (i_icb_rsp_rdata               [  63:   0]),
  .i_icb_rsp_usr                  (i_icb_rsp_usr                 [   2:   0]),
      .o_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .o_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .o_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .o_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .o_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .o_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .o_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .o_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .o_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .o_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .o_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .o_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .o_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .o_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .o_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .o_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .o_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .o_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .o_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .o_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .o_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .o_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .o_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
    wire                splt_bus_icb_cmd_valid        ;
  wire                splt_bus_icb_cmd_ready        ;
  wire                splt_bus_icb_cmd_sel          ;
  wire                splt_bus_icb_cmd_read         ;
  wire    [  31:   0] splt_bus_icb_cmd_addr         ;
  wire    [  63:   0] splt_bus_icb_cmd_wdata        ;
  wire    [   7:   0] splt_bus_icb_cmd_wmask        ;
  wire    [   2:   0] splt_bus_icb_cmd_size         ;
  wire                splt_bus_icb_cmd_lock         ;
  wire                splt_bus_icb_cmd_excl         ;
  wire    [   7:   0] splt_bus_icb_cmd_xlen         ;
  wire    [   1:   0] splt_bus_icb_cmd_xburst       ;
  wire    [   1:   0] splt_bus_icb_cmd_modes        ;
  wire                splt_bus_icb_cmd_dmode        ;
  wire    [   2:   0] splt_bus_icb_cmd_attri        ;
  wire    [   1:   0] splt_bus_icb_cmd_beat         ;
  wire    [   2:   0] splt_bus_icb_cmd_usr          ;
  wire                splt_bus_icb_rsp_ready        ;
  wire                splt_bus_icb_rsp_valid        ;
  wire                splt_bus_icb_rsp_err          ;
  wire                splt_bus_icb_rsp_excl_ok      ;
  wire    [  63:   0] splt_bus_icb_rsp_rdata        ;
  wire    [   2:   0] splt_bus_icb_rsp_usr          ;
      assign                 { o0_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
      assign                 { o0_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
      assign                 { o0_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
      assign                 { o0_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
      assign                 { o0_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
      assign                 { o0_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
      assign                 { o0_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
      assign                 { o0_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
      assign                 { o0_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
      assign                 { o0_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
      assign                 { o0_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
      assign                 { o0_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
      assign                 { o0_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
      assign                 { o0_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
      assign                 { o0_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
      assign                 { o0_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
    assign splt_bus_icb_cmd_ready =
                           { o0_icb_cmd_ready
                           };
    assign splt_bus_icb_rsp_valid =
                           { o0_icb_rsp_valid
                           };
    assign splt_bus_icb_rsp_err =
                           { o0_icb_rsp_err
                           };
    assign splt_bus_icb_rsp_excl_ok =
                           { o0_icb_rsp_excl_ok
                           };
    assign splt_bus_icb_rsp_rdata =
                           { o0_icb_rsp_rdata
                           };
    assign splt_bus_icb_rsp_usr =
                           { o0_icb_rsp_usr
                           };
      assign                 { o0_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
      wire icb_cmd_o0 = 1'b1
                        ; 
  wire [1-1:0] buf_icb_splt_indic = 
      {
                      icb_cmd_o0
      };
  e603_subsys_gnrl_ficb_splt # (
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (SPLT_FIFO_OUTS_NUM ),
  .FIFO_CUT_READY  (SPLT_FIFO_CUT_READY),
  .SPLT_NUM   (1),
  .SPLT_PTR_W (1),
  .SPLT_PTR_1HOT (1),
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .CMD_UW (3),
  .RSP_UW (3),
  .AW         (32),
  .DW         (64) 
  ) u_buf_icb_splt(
      .clk_en(o_clk_en),
  .i_icb_splt_indic       (buf_icb_splt_indic),        
  .splt_active            (splt_active),
      .i_icb_cmd_valid                (buf_icb_cmd_valid                        ),
  .i_icb_cmd_ready                (buf_icb_cmd_ready                        ),
  .i_icb_cmd_sel                  (buf_icb_cmd_sel                          ),
  .i_icb_cmd_read                 (buf_icb_cmd_read                         ),
  .i_icb_cmd_addr                 (buf_icb_cmd_addr              [  31:   0]),
  .i_icb_cmd_wdata                (buf_icb_cmd_wdata             [  63:   0]),
  .i_icb_cmd_wmask                (buf_icb_cmd_wmask             [   7:   0]),
  .i_icb_cmd_size                 (buf_icb_cmd_size              [   2:   0]),
  .i_icb_cmd_lock                 (buf_icb_cmd_lock                         ),
  .i_icb_cmd_excl                 (buf_icb_cmd_excl                         ),
  .i_icb_cmd_xlen                 (buf_icb_cmd_xlen              [   7:   0]),
  .i_icb_cmd_xburst               (buf_icb_cmd_xburst            [   1:   0]),
  .i_icb_cmd_modes                (buf_icb_cmd_modes             [   1:   0]),
  .i_icb_cmd_dmode                (buf_icb_cmd_dmode                        ),
  .i_icb_cmd_attri                (buf_icb_cmd_attri             [   2:   0]),
  .i_icb_cmd_beat                 (buf_icb_cmd_beat              [   1:   0]),
  .i_icb_cmd_usr                  (buf_icb_cmd_usr               [   2:   0]),
  .i_icb_rsp_ready                (buf_icb_rsp_ready                        ),
  .i_icb_rsp_valid                (buf_icb_rsp_valid                        ),
  .i_icb_rsp_err                  (buf_icb_rsp_err                          ),
  .i_icb_rsp_excl_ok              (buf_icb_rsp_excl_ok                      ),
  .i_icb_rsp_rdata                (buf_icb_rsp_rdata             [  63:   0]),
  .i_icb_rsp_usr                  (buf_icb_rsp_usr               [   2:   0]),
      .o_bus_icb_cmd_valid            (splt_bus_icb_cmd_valid                   ),
  .o_bus_icb_cmd_ready            (splt_bus_icb_cmd_ready                   ),
  .o_bus_icb_cmd_sel              (splt_bus_icb_cmd_sel                     ),
  .o_bus_icb_cmd_read             (splt_bus_icb_cmd_read                    ),
  .o_bus_icb_cmd_addr             (splt_bus_icb_cmd_addr         [  31:   0]),
  .o_bus_icb_cmd_wdata            (splt_bus_icb_cmd_wdata        [  63:   0]),
  .o_bus_icb_cmd_wmask            (splt_bus_icb_cmd_wmask        [   7:   0]),
  .o_bus_icb_cmd_size             (splt_bus_icb_cmd_size         [   2:   0]),
  .o_bus_icb_cmd_lock             (splt_bus_icb_cmd_lock                    ),
  .o_bus_icb_cmd_excl             (splt_bus_icb_cmd_excl                    ),
  .o_bus_icb_cmd_xlen             (splt_bus_icb_cmd_xlen         [   7:   0]),
  .o_bus_icb_cmd_xburst           (splt_bus_icb_cmd_xburst       [   1:   0]),
  .o_bus_icb_cmd_modes            (splt_bus_icb_cmd_modes        [   1:   0]),
  .o_bus_icb_cmd_dmode            (splt_bus_icb_cmd_dmode                   ),
  .o_bus_icb_cmd_attri            (splt_bus_icb_cmd_attri        [   2:   0]),
  .o_bus_icb_cmd_beat             (splt_bus_icb_cmd_beat         [   1:   0]),
  .o_bus_icb_cmd_usr              (splt_bus_icb_cmd_usr          [   2:   0]),
  .o_bus_icb_rsp_ready            (splt_bus_icb_rsp_ready                   ),
  .o_bus_icb_rsp_valid            (splt_bus_icb_rsp_valid                   ),
  .o_bus_icb_rsp_err              (splt_bus_icb_rsp_err                     ),
  .o_bus_icb_rsp_excl_ok          (splt_bus_icb_rsp_excl_ok                 ),
  .o_bus_icb_rsp_rdata            (splt_bus_icb_rsp_rdata        [  63:   0]),
  .o_bus_icb_rsp_usr              (splt_bus_icb_rsp_usr          [   2:   0]),
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
`include "global.v"
module e603_subsys_gnrl_rbin4 # (
    parameter ARBT_NUM = 4
)(
  output[ARBT_NUM-1:0] grt_vec,  
  input [ARBT_NUM-1:0] req_vec,  
  input arbt_ena,   
  output rbin4_active,
  input clk,        
  input rst_n
);
  wire [ARBT_NUM-1:0] req_vec_mask;
  wire [ARBT_NUM-1:0] mask_r;
  genvar i;
  generate
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign grt_vec[i] =  ~req_vec_mask[0];
        end
        else if(i==(ARBT_NUM-1)) begin: gen_i_is_msb
          assign grt_vec[i] =  (~(|req_vec[i-1:0])) | req_vec_mask[0];
        end
        else begin:gen_i_is_not_0_and_msb
          assign grt_vec[i] =  (~(|req_vec[i-1:0])) & (~req_vec_mask[i]);
        end
      end
  endgenerate
  localparam CNT_W = 1;
  localparam CNT_1 = 1;
  wire cnt_inc = req_vec[ARBT_NUM-1] & (~grt_vec[ARBT_NUM-1]);
  wire cnt_clr_raw =  grt_vec[ARBT_NUM-1];
  wire mask_set = cnt_inc;
  wire mask_clr = (|mask_r) & cnt_clr_raw;
  wire mask_ena = mask_set | mask_clr;
  wire [ARBT_NUM-1:0] mask_nxt = mask_set ? {1'b0,{ARBT_NUM-1{1'b1}}} : {ARBT_NUM{1'b0}};
e603_subsys_gnrl_dfflr #(ARBT_NUM) mask_dfflr (mask_ena, mask_nxt, mask_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign req_vec_mask = mask_r;
  assign rbin4_active = |mask_r; 
endmodule
`include "global.v"
module e603_subsys_gnrl_ficb_arbt # (
  parameter SUPPORT_LOCK = 1,
  parameter PAYLOAD_NORST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter ARBT_SCHEME = 3,
  parameter RRBIN_CUT_TIMING = 0,
  parameter FIFO_OUTS_NUM = 1,
  parameter FIFO_REG_OUT = 0,
  parameter FIFO_CUT_READY = 0,
  parameter ARBT_NUM = 4,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter ARBT_PTR_W = 2
) (
  output             arbt_active,
  input              clk_en,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [DW-1:0]    o_icb_cmd_wdata,
  output [DW/8-1:0]    o_icb_cmd_wmask,
  output [2-1:0]     o_icb_cmd_beat,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [CMD_SIZE_W-1:0]       o_icb_cmd_size,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  output [ARBT_NUM*1-1:0]     i_bus_icb_cmd_ready,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_valid,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_read,
  input  [ARBT_NUM*AW-1:0]    i_bus_icb_cmd_addr,
  input  [ARBT_NUM*DW-1:0]    i_bus_icb_cmd_wdata,
  input  [ARBT_NUM*DW/8-1:0]    i_bus_icb_cmd_wmask,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_beat ,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_lock ,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_excl ,
  input  [ARBT_NUM*CMD_SIZE_W-1:0]     i_bus_icb_cmd_size ,
  input  [ARBT_NUM*CMD_UW-1:0] i_bus_icb_cmd_usr  ,
  input  [ARBT_NUM*8-1:0]     i_bus_icb_cmd_xlen,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_xburst,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_modes,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_dmode,
  input  [ARBT_NUM*3-1:0]     i_bus_icb_cmd_attri,
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_valid,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_rsp_ready,
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_err,
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_excl_ok,
  output [ARBT_NUM*DW-1:0]    i_bus_icb_rsp_rdata,
  output [ARBT_NUM*RSP_UW-1:0] i_bus_icb_rsp_usr,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_sel_vec,
  input  clk,
  input  rst_n
  );
  localparam ARBT_SCHEME_PRIORITY  = 0;
  localparam ARBT_SCHEME_RROBIN    = 1;
  localparam ARBT_SCHEME_DIRECT_SEL_1HOT = 2;
  localparam ARBT_SCHEME_DIRECT_SEL_PRIORITY = 3;
  localparam ARBT_SCHEME_RROBIN4   = 4;
  localparam ARBT_SCHEME_RROBIN_TIME = 5;
  wire             icb_rsp_valid;
  wire             icb_rsp_ready;
  wire             icb_rsp_err;
  wire             icb_rsp_excl_ok;
  wire [DW-1:0]    icb_rsp_rdata;
  wire [RSP_UW-1:0] icb_rsp_usr;
  wire [ARBT_PTR_W-1:0] t_icb_rsp_id;
  wire                  t_icb_rsp_last;
  localparam RSP_PACK_W = (2+DW+RSP_UW);
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata,
                                 o_icb_rsp_usr};
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 icb_rsp_err,
                                 icb_rsp_excl_ok,
                                 icb_rsp_rdata,
                                 icb_rsp_usr} = rsp_fifo_o_dat;
      assign rsp_fifo_o_dat = rsp_fifo_i_dat;
      assign icb_rsp_valid = o_icb_rsp_valid;
      assign o_icb_rsp_ready = icb_rsp_ready;
  wire rspid_fifo_empty;
  wire rrobin_active;
  wire rrobin_notime_active;
  wire rrobin_time_active;
  wire rbin4_active;
  wire [ARBT_NUM-1:0] lock_mask_r  ;
  wire [ARBT_NUM-1:0] omask_r;
  wire [ARBT_NUM-1:0] burst_mask_r;
genvar i;
generate 
  if(ARBT_NUM == 1) begin:gen_arbt_num_eq_1
    assign i_bus_icb_cmd_ready = o_icb_cmd_ready    ;
    assign o_icb_cmd_valid     = i_bus_icb_cmd_valid;
    assign o_icb_cmd_sel       = i_bus_icb_cmd_sel_vec  ;
    assign o_icb_cmd_read      = i_bus_icb_cmd_read ;
    assign o_icb_cmd_addr      = i_bus_icb_cmd_addr ;
    assign o_icb_cmd_wdata     = i_bus_icb_cmd_wdata;
    assign o_icb_cmd_wmask     = i_bus_icb_cmd_wmask;
    assign o_icb_cmd_beat      = i_bus_icb_cmd_beat ;
    assign o_icb_cmd_lock      = i_bus_icb_cmd_lock ;
    assign o_icb_cmd_excl      = i_bus_icb_cmd_excl ;
    assign o_icb_cmd_size      = i_bus_icb_cmd_size ;
    assign o_icb_cmd_usr       = i_bus_icb_cmd_usr  ;
    assign o_icb_cmd_xlen      = i_bus_icb_cmd_xlen  ;
    assign o_icb_cmd_xburst    = i_bus_icb_cmd_xburst;
    assign o_icb_cmd_modes     = i_bus_icb_cmd_modes ;
    assign o_icb_cmd_dmode     = i_bus_icb_cmd_dmode ;
    assign o_icb_cmd_attri     = i_bus_icb_cmd_attri ;
    assign icb_rsp_ready     = i_bus_icb_rsp_ready;
    assign i_bus_icb_rsp_valid = icb_rsp_valid    ;
    assign i_bus_icb_rsp_err   = icb_rsp_err      ;
    assign i_bus_icb_rsp_excl_ok   = icb_rsp_excl_ok      ;
    assign i_bus_icb_rsp_rdata = icb_rsp_rdata    ;
    assign i_bus_icb_rsp_usr   = icb_rsp_usr      ;
    assign rspid_fifo_empty    = 1'b1;
    assign lock_mask_r = {ARBT_NUM{1'b0}};
    assign omask_r = {ARBT_NUM{1'b0}};
    assign burst_mask_r = {ARBT_NUM{1'b0}};
    assign rbin4_active = 1'b0;
    assign rrobin_active = 1'b0;
    assign rrobin_time_active = 1'b0;
    assign rrobin_notime_active = 1'b0;
  end
  else begin:gen_arbt_num_gt_1
    integer j;
    wire [ARBT_NUM-1:0] i_bus_icb_cmd_grt_vec;
    wire [ARBT_NUM-1:0] i_bus_icb_cmd_sel;
    wire o_icb_cmd_valid_real;
    wire o_icb_cmd_ready_real;
    wire            i_icb_cmd_read [ARBT_NUM-1:0];
    wire [AW-1:0]   i_icb_cmd_addr [ARBT_NUM-1:0];
    wire [DW-1:0]   i_icb_cmd_wdata[ARBT_NUM-1:0];
    wire [DW/8-1:0]   i_icb_cmd_wmask[ARBT_NUM-1:0];
    wire [2-1:0]    i_icb_cmd_beat [ARBT_NUM-1:0];
    wire            i_icb_cmd_lock [ARBT_NUM-1:0];
    wire            i_icb_cmd_excl [ARBT_NUM-1:0];
    wire [CMD_SIZE_W-1:0]    i_icb_cmd_size [ARBT_NUM-1:0];
    wire [CMD_UW-1:0]i_icb_cmd_usr  [ARBT_NUM-1:0];
    wire [7:0]      i_icb_cmd_xlen   [ARBT_NUM-1:0];
    wire [1:0]      i_icb_cmd_xburst [ARBT_NUM-1:0];
    wire [1:0]      i_icb_cmd_modes  [ARBT_NUM-1:0];
    wire            i_icb_cmd_dmode  [ARBT_NUM-1:0];
    wire [2:0]      i_icb_cmd_attri  [ARBT_NUM-1:0];
    reg            sel_o_icb_cmd_read;
    reg [AW-1:0]   sel_o_icb_cmd_addr;
    reg [DW-1:0]   sel_o_icb_cmd_wdata;
    reg [DW/8-1:0]   sel_o_icb_cmd_wmask;
    reg [2-1:0]    sel_o_icb_cmd_beat ;
    reg            sel_o_icb_cmd_lock ;
    reg            sel_o_icb_cmd_excl ;
    reg [CMD_SIZE_W-1:0]    sel_o_icb_cmd_size ;
    reg [CMD_UW-1:0]sel_o_icb_cmd_usr  ;
    reg [7:0]      sel_o_icb_cmd_xlen  ;
    reg [1:0]      sel_o_icb_cmd_xburst;
    reg [1:0]      sel_o_icb_cmd_modes ;
    reg            sel_o_icb_cmd_dmode ;
    reg [2:0]      sel_o_icb_cmd_attri ;
    wire icb_rsp_ready_pre;
    wire icb_rsp_valid_pre;
    wire rspid_fifo_bypass;
    wire rspid_fifo_wen;
    wire rspid_fifo_ren;
    wire rspid_fifo_i_valid;
    wire rspid_fifo_o_valid;
    wire rspid_fifo_i_ready;
    wire rspid_fifo_o_ready;
    wire [ARBT_PTR_W-1:0] rspid_fifo_rdat;
    wire [ARBT_PTR_W-1:0] rspid_fifo_wdat;
    wire rspid_fifo_full;
    reg [ARBT_PTR_W-1:0] i_arbt_indic_id;
    wire [ARBT_NUM*1-1:0] i_bus_icb_cmd_ready_pos;
    wire [ARBT_NUM*1-1:0] i_bus_icb_cmd_valid_pos;
    wire [ARBT_NUM*1-1:0] i_bus_icb_cmd_sel_vec_pos;
    wire arbt_ena;
    wire [ARBT_PTR_W-1:0] icb_rsp_port_id;
    if((ARBT_SCHEME == ARBT_SCHEME_RROBIN) || (ARBT_SCHEME == ARBT_SCHEME_RROBIN_TIME) || (ARBT_SCHEME == ARBT_SCHEME_RROBIN4)) begin: gen_rrobin
        assign omask_r = {ARBT_NUM{1'b0}};
    end
    else begin: gen_not_rrobin
        wire [ARBT_NUM-1:0] omask_nxt;
        wire omask_ena;
        wire omask_set;
        wire omask_clr;
        assign omask_set = o_icb_cmd_valid_real & (~arbt_ena); 
        assign omask_clr = (|omask_r) & (arbt_ena | (~o_icb_cmd_valid_real));
        assign omask_ena = clk_en & (omask_set | omask_clr);
        assign omask_nxt = omask_clr ? {ARBT_NUM{1'b0}} : (~i_bus_icb_cmd_sel); 
e603_subsys_gnrl_dfflr #(ARBT_NUM) omask_dfflr (omask_ena, omask_nxt, omask_r, clk, rst_n);// VPP_NO_REG_PARSE
    end
    wire [ARBT_NUM-1:0] burst_mask_nxt;
    wire burst_mask_ena;
    wire burst_mask_set;
    wire burst_mask_clr;
      assign burst_mask_set = o_icb_cmd_beat[0] & arbt_ena;
      assign burst_mask_clr = (|burst_mask_r) & o_icb_cmd_beat[1] & arbt_ena;
    assign burst_mask_ena = clk_en & (burst_mask_set | burst_mask_clr);
    assign burst_mask_nxt = burst_mask_clr ? {ARBT_NUM{1'b0}} : (~i_bus_icb_cmd_sel); 
e603_subsys_gnrl_dfflr #(ARBT_NUM) burst_mask_dfflr (burst_mask_ena, burst_mask_nxt, burst_mask_r, clk, rst_n);// VPP_NO_REG_PARSE
      assign i_bus_icb_cmd_valid_pos   = (~burst_mask_r) & (~omask_r) & (~lock_mask_r) & i_bus_icb_cmd_valid;
      assign i_bus_icb_cmd_ready       = (~burst_mask_r) & (~omask_r) & (~lock_mask_r) & i_bus_icb_cmd_ready_pos;
      assign i_bus_icb_cmd_sel_vec_pos = (~burst_mask_r) & (~omask_r) & (~lock_mask_r) & i_bus_icb_cmd_sel_vec;
    assign o_icb_cmd_sel   = |i_bus_icb_cmd_sel_vec_pos;
    assign o_icb_cmd_valid = o_icb_cmd_valid_real & (~rspid_fifo_full);
    assign o_icb_cmd_ready_real = o_icb_cmd_ready & (~rspid_fifo_full);
    for(i = 0; i < ARBT_NUM; i = i+1)
    begin:gen_icb_distract
      assign i_icb_cmd_read [i] = i_bus_icb_cmd_read [(i+1)*1     -1 : i*1     ];
      assign i_icb_cmd_addr [i] = i_bus_icb_cmd_addr [(i+1)*AW    -1 : i*AW    ];
      assign i_icb_cmd_wdata[i] = i_bus_icb_cmd_wdata[(i+1)*DW    -1 : i*DW    ];
      assign i_icb_cmd_wmask[i] = i_bus_icb_cmd_wmask[(i+1)*DW/8    -1 : i*DW/8    ];
      assign i_icb_cmd_beat [i] = i_bus_icb_cmd_beat [(i+1)*2     -1 : i*2     ];
      assign i_icb_cmd_lock [i] = i_bus_icb_cmd_lock [(i+1)*1     -1 : i*1     ];
      assign i_icb_cmd_excl [i] = i_bus_icb_cmd_excl [(i+1)*1     -1 : i*1     ];
      assign i_icb_cmd_size [i] = i_bus_icb_cmd_size [(i+1)*CMD_SIZE_W     -1 : i*CMD_SIZE_W     ];
      assign i_icb_cmd_usr  [i] = i_bus_icb_cmd_usr  [(i+1)*CMD_UW -1 : i*CMD_UW ];
      assign i_icb_cmd_xlen  [i] = i_bus_icb_cmd_xlen   [(i+1)*8 -1 : i*8 ];
      assign i_icb_cmd_xburst[i] = i_bus_icb_cmd_xburst [(i+1)*2 -1 : i*2 ];
      assign i_icb_cmd_modes [i] = i_bus_icb_cmd_modes  [(i+1)*2 -1 : i*2 ];
      assign i_icb_cmd_dmode [i] = i_bus_icb_cmd_dmode  [(i+1)*1 -1 : i*1 ];
      assign i_icb_cmd_attri [i] = i_bus_icb_cmd_attri  [(i+1)*3 -1 : i*3 ];
      assign i_bus_icb_cmd_ready_pos[i] = i_bus_icb_cmd_grt_vec[i] & o_icb_cmd_ready_real;
      assign i_bus_icb_rsp_valid[i] = icb_rsp_valid_pre & (icb_rsp_port_id == i[ARBT_PTR_W-1:0]);
    end
    assign arbt_ena = o_icb_cmd_valid & o_icb_cmd_ready;
      wire [ARBT_NUM-1:0] lock_mask_set;
      wire [ARBT_NUM-1:0] lock_mask_clr;
      wire [ARBT_NUM-1:0] lock_mask_ena;
      wire [ARBT_NUM-1:0] lock_mask_nxt;
      for(i = 0; i < ARBT_NUM; i = i+1) begin:gen_lock_mask
        assign lock_mask_set[i] = clk_en & (i_bus_icb_cmd_sel[i] == 1'b0) & o_icb_cmd_lock & arbt_ena;
        assign lock_mask_clr[i] = clk_en & lock_mask_r[i] & ((~o_icb_cmd_lock) & arbt_ena);
        assign lock_mask_ena[i] = lock_mask_set[i] |   lock_mask_clr[i];
        assign lock_mask_nxt[i] = lock_mask_set[i] & (~lock_mask_clr[i]);
        if(SUPPORT_LOCK == 1) begin: support_lock_gen
e603_subsys_gnrl_dfflr #(1) lock_mask_dfflr (lock_mask_ena[i], lock_mask_nxt[i], lock_mask_r[i], clk, rst_n);// VPP_NO_REG_PARSE
        end
        else begin: no_support_lock_gen
        assign lock_mask_r[i] = 1'b0;
        end
      end
    if(ARBT_SCHEME == ARBT_SCHEME_PRIORITY) begin:gen_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_icb_cmd_grt_vec[i] =  1'b1;
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_valid_pos[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_icb_cmd_grt_vec[i] =  ~(|i_bus_icb_cmd_valid_pos[i-1:0]);
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_valid_pos[i];
        end
      end
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN) begin:gen_rrobin_arbt
       if(RRBIN_CUT_TIMING == 1) begin:gen_rbin_cut_timing
      wire lock_mask_r_set  = |(lock_mask_set & (~lock_mask_clr));
      wire burst_mask_r_set = |(burst_mask_set & (~burst_mask_clr));
     e603_subsys_gnrl_rrobin_cut # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin_cut(
       .rrobin_active (rrobin_notime_active),
       .grt_vec  (i_bus_icb_cmd_grt_vec),
       .req_vec  (i_bus_icb_cmd_sel_vec_pos),
       .req_mask  (burst_mask_r | lock_mask_r),
       .req_mask_set  (burst_mask_r_set | lock_mask_r_set),
       .arbt_ena (arbt_ena & clk_en),
       .clk      (clk),
       .rst_n    (rst_n)
     );
       end
       else begin: no_gen_rbin_cut_ciming
     e603_subsys_gnrl_rrobin # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin(
       .rrobin_active (rrobin_notime_active),
       .grt_vec  (i_bus_icb_cmd_grt_vec),
       .req_vec  (i_bus_icb_cmd_sel_vec_pos),
       .arbt_ena (arbt_ena & clk_en),
       .clk      (clk),
       .rst_n    (rst_n)
     );
       end
     assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec;
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
   end
   else begin: gen_no_rrobin
     assign rrobin_notime_active = 1'b0;
   end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN_TIME) begin:gen_rrobin_time_arbt
     e603_subsys_gnrl_rrobin_time # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin_time(
       .rrobin_active (rrobin_time_active),
       .grt_vec  (i_bus_icb_cmd_grt_vec),
       .req_vec  (i_bus_icb_cmd_valid),
       .req_mask  (burst_mask_r | lock_mask_r),
       .arbt_ena (arbt_ena & clk_en),
       .clk      (clk),
       .rst_n    (rst_n)
     );
     assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec;
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid & i_bus_icb_cmd_sel);
   end
   else begin: gen_no_rrobin_time
     assign rrobin_time_active = 1'b0;
   end
   assign rrobin_active = rrobin_notime_active | rrobin_time_active | rbin4_active;
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_1HOT) begin:gen_indic_arbt
     assign i_bus_icb_cmd_grt_vec = i_bus_icb_cmd_sel_vec_pos;
     assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec;
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
   end
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_PRIORITY) begin:gen_indic_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_icb_cmd_grt_vec[i] =  1'b1;
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_sel_vec_pos[i];
        end
        else if(i==(ARBT_NUM-1)) begin: gen_i_is_n
          assign i_bus_icb_cmd_grt_vec[i] =  ~(|i_bus_icb_cmd_sel_vec_pos[i-1:0]);
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_icb_cmd_grt_vec[i] =  ~(|i_bus_icb_cmd_sel_vec_pos[i-1:0]);
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_sel_vec_pos[i];
        end
      end
      assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN4) begin:gen_rbin4_arbt
      wire lock_mask_r_set  = |lock_mask_set ;
      wire burst_mask_r_set = |burst_mask_set;
      e603_subsys_gnrl_rbin4 # (
          .ARBT_NUM(ARBT_NUM)
      )u_e603_subsys_gnrl_rbin4(
        .grt_vec  (i_bus_icb_cmd_grt_vec),
        .req_vec  (i_bus_icb_cmd_sel_vec_pos),
        .arbt_ena (arbt_ena & clk_en & (~lock_mask_r_set) & (~burst_mask_r_set)),
        .rbin4_active(rbin4_active),
        .clk      (clk),
        .rst_n    (rst_n)
      );
      assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec & i_bus_icb_cmd_sel_vec_pos;
      assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
   end
   else begin:gen_no_rbin4_arbt
      assign rbin4_active = 1'b0;
   end
    always @ (*) begin : sel_o_icb_cmd_ready_PROC
      sel_o_icb_cmd_read  = {1   {1'b0}};
      sel_o_icb_cmd_addr  = {AW  {1'b0}};
      sel_o_icb_cmd_wdata = {DW  {1'b0}};
      sel_o_icb_cmd_wmask = {DW/8  {1'b0}};
      sel_o_icb_cmd_beat  = {2   {1'b0}};
      sel_o_icb_cmd_lock  = {1   {1'b0}};
      sel_o_icb_cmd_excl  = {1   {1'b0}};
      sel_o_icb_cmd_size  = {CMD_SIZE_W   {1'b0}};
      sel_o_icb_cmd_usr   = {CMD_UW{1'b0}};
      sel_o_icb_cmd_xlen  = {8{1'b0}};
      sel_o_icb_cmd_xburst= {2{1'b0}};
      sel_o_icb_cmd_modes = {2{1'b0}};
      sel_o_icb_cmd_dmode = {1{1'b0}};
      sel_o_icb_cmd_attri = {3{1'b0}};
      for(j = 0; j < ARBT_NUM; j = j+1) begin
        sel_o_icb_cmd_read  = sel_o_icb_cmd_read  | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_read [j]);
        sel_o_icb_cmd_addr  = sel_o_icb_cmd_addr  | ({AW   {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_addr [j]);
        sel_o_icb_cmd_wdata = sel_o_icb_cmd_wdata | ({DW   {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_wdata[j]);
        sel_o_icb_cmd_wmask = sel_o_icb_cmd_wmask | ({DW/8   {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_wmask[j]);
        sel_o_icb_cmd_beat  = sel_o_icb_cmd_beat  | ({2    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_beat [j]);
        sel_o_icb_cmd_lock  = sel_o_icb_cmd_lock  | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_lock [j]);
        sel_o_icb_cmd_excl  = sel_o_icb_cmd_excl  | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_excl [j]);
        sel_o_icb_cmd_size  = sel_o_icb_cmd_size  | ({CMD_SIZE_W    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_size [j]);
        sel_o_icb_cmd_usr   = sel_o_icb_cmd_usr   | ({CMD_UW{i_bus_icb_cmd_sel[j]}} & i_icb_cmd_usr  [j]);
        sel_o_icb_cmd_xlen  = sel_o_icb_cmd_xlen  | ({8    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_xlen  [j]);
        sel_o_icb_cmd_xburst= sel_o_icb_cmd_xburst| ({2    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_xburst[j]);
        sel_o_icb_cmd_modes = sel_o_icb_cmd_modes | ({2    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_modes [j]);
        sel_o_icb_cmd_dmode = sel_o_icb_cmd_dmode | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_dmode [j]);
        sel_o_icb_cmd_attri = sel_o_icb_cmd_attri | ({3    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_attri [j]);
      end
    end
    always @ (*) begin : i_arbt_indic_id_PROC
      i_arbt_indic_id = {ARBT_PTR_W{1'b0}};
      for(j = 0; j < ARBT_NUM; j = j+1) begin
// spyglass disable_block W216
// SMD: Inappropriate range select for int_part_sel variable
// SJ:  Here is not a real issue
        i_arbt_indic_id = i_arbt_indic_id | ({ARBT_PTR_W{i_bus_icb_cmd_sel[j]}} & (j[ARBT_PTR_W-1:0]));
// spyglass enable_block W216
      end
    end
    assign rspid_fifo_wen = o_icb_cmd_valid & o_icb_cmd_ready;
    assign rspid_fifo_ren = icb_rsp_valid & icb_rsp_ready;
    if(ALLOW_0CYCL_RSP == 1) begin: gen_allow_0rsp
        assign rspid_fifo_bypass = rspid_fifo_empty & rspid_fifo_wen & rspid_fifo_ren;
        assign icb_rsp_port_id = rspid_fifo_empty ? rspid_fifo_wdat : rspid_fifo_rdat;
        assign icb_rsp_valid_pre = icb_rsp_valid;
        assign icb_rsp_ready     = icb_rsp_ready_pre;
    end
    else begin: gen_no_allow_0rsp
        assign rspid_fifo_bypass   = 1'b0;
        assign icb_rsp_port_id   = rspid_fifo_rdat;
        assign icb_rsp_valid_pre = (~rspid_fifo_empty) & icb_rsp_valid;
        assign icb_rsp_ready     = (~rspid_fifo_empty) & icb_rsp_ready_pre;
    end
    assign rspid_fifo_i_valid = clk_en & rspid_fifo_wen & (~rspid_fifo_bypass);
    assign rspid_fifo_full    = (~rspid_fifo_i_ready);
    assign rspid_fifo_o_ready = clk_en & rspid_fifo_ren & (~rspid_fifo_bypass);
    assign rspid_fifo_empty   = (~rspid_fifo_o_valid);
    assign rspid_fifo_wdat   = i_arbt_indic_id;
    if(FIFO_OUTS_NUM == 1) begin:gen_dp_1
      e603_subsys_gnrl_pipe_stage # (
        .CUT_READY (FIFO_CUT_READY),
        .DP  (1),
        .DW  (ARBT_PTR_W)
      ) u_e603_subsys_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else begin: gen_dp_gt1
      e603_subsys_gnrl_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT(FIFO_REG_OUT),
        .CUT_READY(FIFO_CUT_READY),
        .DP  (FIFO_OUTS_NUM),
        .DW  (ARBT_PTR_W)
      ) u_e603_subsys_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    assign o_icb_cmd_read  = sel_o_icb_cmd_read ;
    assign o_icb_cmd_addr  = sel_o_icb_cmd_addr ;
    assign o_icb_cmd_wdata = sel_o_icb_cmd_wdata;
    assign o_icb_cmd_wmask = sel_o_icb_cmd_wmask;
    assign o_icb_cmd_beat  = sel_o_icb_cmd_beat ;
    assign o_icb_cmd_lock  = sel_o_icb_cmd_lock ;
    assign o_icb_cmd_excl  = sel_o_icb_cmd_excl ;
    assign o_icb_cmd_size  = sel_o_icb_cmd_size ;
    assign o_icb_cmd_usr   = sel_o_icb_cmd_usr  ;
    assign o_icb_cmd_xlen  = sel_o_icb_cmd_xlen  ;
    assign o_icb_cmd_xburst= sel_o_icb_cmd_xburst;
    assign o_icb_cmd_modes = sel_o_icb_cmd_modes ;
    assign o_icb_cmd_dmode = sel_o_icb_cmd_dmode ;
    assign o_icb_cmd_attri = sel_o_icb_cmd_attri ;
    assign icb_rsp_ready_pre = i_bus_icb_rsp_ready[icb_rsp_port_id];
    assign i_bus_icb_rsp_err     = {ARBT_NUM{icb_rsp_err  }};
    assign i_bus_icb_rsp_excl_ok = {ARBT_NUM{icb_rsp_excl_ok}};
    assign i_bus_icb_rsp_rdata   = {ARBT_NUM{icb_rsp_rdata}};
    assign i_bus_icb_rsp_usr     = {ARBT_NUM{icb_rsp_usr}};
  end
  endgenerate 
  assign arbt_active =
         (|i_bus_icb_cmd_sel_vec) | (~rspid_fifo_empty) | icb_rsp_valid | (|burst_mask_r)| (|omask_r) | (|lock_mask_r) | rrobin_active;
endmodule
module e603_subsys_gnrl_ficb_buffer # (
    parameter OUTS_CNT_BLOCK_THROUGH = 0,
    parameter RSP_STRICT_ORDER = 0,
  parameter PAYLOAD_NORST = 0,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter CMD_MSKO = 0,
  parameter OUTS_CNT_W = 1,
  parameter AW = 32,
  parameter DW = 32,
  parameter CMD_CUT_READY = 0,
  parameter RSP_CUT_READY = 0,
  parameter ACTIVE_USE_FLOP_CLEAN = 0,
  parameter CMD_DP = 0,
  parameter RSP_DP = 0,
  parameter CMD_BYPBUF = 0,
  parameter CMD_RGLR_FIFO = 0,
  parameter RSP_BYPBUF = 0,
  parameter RSP_RGLR_FIFO = 0,
  parameter REG_OUT = 0,
  parameter RSP_ALWAYS_READY = 0,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  input              i_clk_en,
  input              o_clk_en,
  output             icb_buffer_active,
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [DW-1:0]    i_icb_cmd_wdata,
  input  [DW/8-1:0]  i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [DW-1:0]    i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [DW-1:0]    o_icb_cmd_wdata,
  output [DW/8-1:0]  o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  localparam CMD_PACK_W = (1+AW+DW+DW/8+1+3+3+CMD_UW+8+2+2+1+3 + 0);
  localparam RSP_PACK_W = (2+DW+RSP_UW + 0);
 wire i_icb_cmd_xlen_eq0 = (i_icb_cmd_xlen == 8'd0);
 wire i_icb_cmd_first = i_icb_cmd_beat[0] | i_icb_cmd_xlen_eq0;
 wire o_icb_cmd_xlen_eq0 = (o_icb_cmd_xlen == 8'd0);
 wire o_icb_cmd_first = o_icb_cmd_beat[0] | o_icb_cmd_xlen_eq0;
 generate
   if((CMD_DP == 0) && (RSP_DP == 0)) begin:gen_icb_buf_through
  wire outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready & i_clk_en 
    ;
  wire outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & i_clk_en 
    ;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
      assign icb_buffer_active =
      i_icb_cmd_sel | (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
    wire i_outs_cnt_is_max;
    if(OUTS_CNT_BLOCK_THROUGH == 1) begin:outs_cnt_block_through
        assign i_outs_cnt_is_max = (outs_cnt_r == {OUTS_CNT_W{1'b1}});
    end
    else begin:outs_cnt_no_block_through
        assign i_outs_cnt_is_max = 1'b0;
    end
    assign i_icb_cmd_ready = (~i_outs_cnt_is_max) & o_icb_cmd_ready;
    assign o_icb_cmd_sel   = (~i_outs_cnt_is_max) & i_icb_cmd_sel;
    assign o_icb_cmd_valid = (~i_outs_cnt_is_max) & i_icb_cmd_valid;
    assign o_icb_cmd_read  = i_icb_cmd_read ;
    assign o_icb_cmd_addr  = i_icb_cmd_addr ;
    assign o_icb_cmd_wdata = i_icb_cmd_wdata;
    assign o_icb_cmd_wmask = i_icb_cmd_wmask;
    assign o_icb_cmd_beat  = i_icb_cmd_beat ;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
    assign o_icb_cmd_size  = o_icb_cmd_size_pre ;
    assign o_icb_cmd_xlen  = o_icb_cmd_xlen_pre  ;
    assign o_icb_cmd_lock  = i_icb_cmd_lock ;
    assign o_icb_cmd_excl  = i_icb_cmd_excl ;
    assign o_icb_cmd_size_pre  = i_icb_cmd_size ;
    assign o_icb_cmd_usr   = i_icb_cmd_usr  ;
    assign o_icb_cmd_xlen_pre  = i_icb_cmd_xlen  ;
    assign o_icb_cmd_xburst= i_icb_cmd_xburst;
    assign o_icb_cmd_modes = i_icb_cmd_modes ;
    assign o_icb_cmd_dmode = i_icb_cmd_dmode ;
    assign o_icb_cmd_attri = i_icb_cmd_attri ;
    assign o_icb_rsp_ready = i_icb_rsp_ready;
    assign i_icb_rsp_valid     = o_icb_rsp_valid;
    assign i_icb_rsp_err       = o_icb_rsp_err  ;
    assign i_icb_rsp_excl_ok   = o_icb_rsp_excl_ok  ;
    assign i_icb_rsp_rdata     = o_icb_rsp_rdata;
    assign i_icb_rsp_usr       = o_icb_rsp_usr;
  end
  else begin:gen_icb_buf_not_through
  wire [CMD_PACK_W-1:0] cmd_fifo_i_dat = {
                                 i_icb_cmd_read,
                                 i_icb_cmd_addr,
                                 i_icb_cmd_wdata,
                                 i_icb_cmd_wmask,
                                 i_icb_cmd_lock,
                                 i_icb_cmd_excl,
                                 i_icb_cmd_size,
                                 i_icb_cmd_beat,
                                 i_icb_cmd_xlen,
                                 i_icb_cmd_xburst,
                                 i_icb_cmd_modes,
                                 i_icb_cmd_dmode,
                                 i_icb_cmd_attri,
                                 i_icb_cmd_usr};
  wire [CMD_PACK_W-1:0] cmd_fifo_o_dat;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
    assign o_icb_cmd_size  = o_icb_cmd_size_pre ;
    assign o_icb_cmd_xlen  = o_icb_cmd_xlen_pre  ;
  assign {
                                 o_icb_cmd_read,
                                 o_icb_cmd_addr,
                                 o_icb_cmd_wdata,
                                 o_icb_cmd_wmask,
                                 o_icb_cmd_lock,
                                 o_icb_cmd_excl,
                                 o_icb_cmd_size_pre,
                                 o_icb_cmd_beat,
                                 o_icb_cmd_xlen_pre,
                                 o_icb_cmd_xburst,
                                 o_icb_cmd_modes,
                                 o_icb_cmd_dmode,
                                 o_icb_cmd_attri,
                                 o_icb_cmd_usr} = cmd_fifo_o_dat;
  wire o_icb_cmd_valid_pre;
  wire o_icb_cmd_ready_pre;
  wire outs_cnt_full;
  wire cmd_fifo_i_valid;
  wire cmd_fifo_i_ready;
  assign cmd_fifo_i_valid = (~outs_cnt_full) & i_icb_cmd_valid;
  assign i_icb_cmd_ready  = (~outs_cnt_full) & cmd_fifo_i_ready;
  wire cmd_ratio_fifo_active;
    if(CMD_RGLR_FIFO == 1) begin: gen_cmd_rlgr_fifo
  e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP  (CMD_DP),
    .DW  (CMD_PACK_W)
  ) u_e603_subsys_gnrl_cmd_fifo (
    .i_vld(cmd_fifo_i_valid),
    .i_rdy(cmd_fifo_i_ready),
    .i_dat(cmd_fifo_i_dat ),
    .o_vld(o_icb_cmd_valid_pre),
    .o_rdy(o_icb_cmd_ready_pre),
    .o_dat(cmd_fifo_o_dat ),
    .clk  (clk),
    .rst_n(rst_n)
  );
   assign cmd_ratio_fifo_active = o_icb_cmd_valid_pre;
    end
    else if(CMD_BYPBUF == 0) begin: gen_cmd_no_bypbuf
  e603_subsys_gnrl_ratio_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .I_SUPPORT_RATIO (I_SUPPORT_RATIO),
        .O_SUPPORT_RATIO (O_SUPPORT_RATIO),
    .DP  (CMD_DP),
    .DW  (CMD_PACK_W)
  ) u_e603_subsys_gnrl_cmd_fifo (
    .i_clk_en     (i_clk_en),
    .o_clk_en     (o_clk_en),
    .o_fifo_active(cmd_ratio_fifo_active),
    .i_vld(cmd_fifo_i_valid),
    .i_rdy(cmd_fifo_i_ready),
    .i_dat(cmd_fifo_i_dat ),
    .o_vld(o_icb_cmd_valid_pre),
    .o_rdy(o_icb_cmd_ready_pre),
    .o_dat(cmd_fifo_o_dat ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    else begin:gen_cmd_bypbuf
  e603_subsys_gnrl_bypbuf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP  (CMD_DP),
    .DW  (CMD_PACK_W)
  ) u_e603_subsys_gnrl_cmd_bypbuf (
    .i_vld(cmd_fifo_i_valid & i_clk_en),
    .i_rdy(cmd_fifo_i_ready),
    .i_dat(cmd_fifo_i_dat ),
    .o_vld(o_icb_cmd_valid_pre),
    .o_rdy(o_icb_cmd_ready_pre & o_clk_en),
    .o_dat(cmd_fifo_o_dat ),
        .fifo_o_vld(cmd_ratio_fifo_active),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
   wire oo_outs_cnt_max;
   wire o_outs_cnt_max;
    if(CMD_DP == 0) begin:dp_is_0_gen
        assign o_icb_cmd_sel = i_icb_cmd_sel;
    end
    else begin:dp_is_not_0_gen
        assign o_icb_cmd_sel = o_icb_cmd_valid_pre;
    end
  wire rsp_buf_ready;
    if(RSP_ALWAYS_READY == 1) begin: gen_rsp_always_ready_1
      assign o_icb_cmd_valid     = rsp_buf_ready & o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = rsp_buf_ready & o_icb_cmd_ready;
    end
    else begin: gen_rsp_always_ready_0
      assign o_icb_cmd_valid     = o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = o_icb_cmd_ready;
    end
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata,
                                 o_icb_rsp_usr};
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 i_icb_rsp_err,
                                 i_icb_rsp_excl_ok,
                                 i_icb_rsp_rdata,
                                 i_icb_rsp_usr} = rsp_fifo_o_dat;
  wire o_icb_rsp_valid_raw;
  wire o_icb_rsp_ready_raw;
    if(RSP_RGLR_FIFO == 1) begin: gen_rsp_rlgr_fifo
      e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT (REG_OUT),
        .DP  (RSP_DP),
        .DW  (RSP_PACK_W)
      ) u_e603_subsys_gnrl_rsp_fifo (
        .i_vld(o_icb_rsp_valid_raw),
        .i_rdy(o_icb_rsp_ready_raw),
        .i_dat(rsp_fifo_i_dat ),
        .o_vld(i_icb_rsp_valid),
        .o_rdy(i_icb_rsp_ready),
        .o_dat(rsp_fifo_o_dat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else if(RSP_BYPBUF == 0) begin: gen_rsp_no_bypbuf
      e603_subsys_gnrl_ratio_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .I_SUPPORT_RATIO (O_SUPPORT_RATIO),
        .O_SUPPORT_RATIO (I_SUPPORT_RATIO),
        .REG_OUT (REG_OUT),
        .DP  (RSP_DP),
        .DW  (RSP_PACK_W)
      ) u_e603_subsys_gnrl_rsp_fifo (
        .i_clk_en     (o_clk_en),
        .o_clk_en     (i_clk_en),
        .o_fifo_active(),
        .i_vld(o_icb_rsp_valid_raw),
        .i_rdy(o_icb_rsp_ready_raw),
        .i_dat(rsp_fifo_i_dat ),
        .o_vld(i_icb_rsp_valid),
        .o_rdy(i_icb_rsp_ready),
        .o_dat(rsp_fifo_o_dat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else begin:gen_rsp_bypbuf
      e603_subsys_gnrl_bypbuf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RSP_DP),
        .DW  (RSP_PACK_W)
      ) u_e603_subsys_gnrl_rsp_bypbuf (
        .i_vld(o_icb_rsp_valid_raw & o_clk_en),
        .i_rdy(o_icb_rsp_ready_raw),
        .i_dat(rsp_fifo_i_dat ),
        .o_vld(i_icb_rsp_valid),
        .o_rdy(i_icb_rsp_ready & i_clk_en),
        .o_dat(rsp_fifo_o_dat ),
        .fifo_o_vld(),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
  wire outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready & i_clk_en
                    ;
  wire outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & i_clk_en
                    ;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign outs_cnt_full = (outs_cnt_r == {OUTS_CNT_W{1'b1}});
   if((CMD_BYPBUF != 1) && (CMD_DP != 0) && (ACTIVE_USE_FLOP_CLEAN == 1)) begin:gen_active_flop_clean
  assign icb_buffer_active =
      (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
   end
   else begin: gen_active_no_flop_clean
  assign icb_buffer_active =
      i_icb_cmd_sel | cmd_ratio_fifo_active | (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
   end
  wire o_outs_cnt_inc = o_icb_cmd_valid & o_icb_cmd_ready & o_clk_en 
                    ;
  wire o_outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & i_clk_en 
                    ;
  wire o_outs_cnt_ena = o_outs_cnt_inc ^ o_outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_r;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_nxt = o_outs_cnt_inc ? (o_outs_cnt_r + 1'b1) : (o_outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) o_outs_cnt_dfflr (o_outs_cnt_ena, o_outs_cnt_nxt, o_outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire [OUTS_CNT_W-1:0] o_outs_cnt_din = o_outs_cnt_ena ? o_outs_cnt_nxt : o_outs_cnt_r;
  wire rsp_buf_ready_raw = ~(o_outs_cnt_r   == RSP_DP[OUTS_CNT_W-1:0]);
  wire rsp_buf_ready_din = ~(o_outs_cnt_din == RSP_DP[OUTS_CNT_W-1:0]);
    wire o_need_updat = o_outs_cnt_ena;
    wire o_need_updat_r;
    wire o_need_updat_r_set = (o_need_updat && !o_clk_en);
    wire o_need_updat_r_clr = (o_need_updat_r && o_clk_en);
    wire o_need_updat_r_ena = o_need_updat_r_set || o_need_updat_r_clr;
    wire o_need_updat_r_nxt = o_need_updat_r_set;
e603_subsys_gnrl_dfflr  #(1) o_need_updat_r_dfflr    (o_need_updat_r_ena, o_need_updat_r_nxt, o_need_updat_r,     clk, rst_n);// VPP_NO_REG_PARSE
    wire rsp_buf_ready_r;
    wire rsp_buf_ready_r_ena = o_clk_en && (o_need_updat || o_need_updat_r);
    wire rsp_buf_ready_r_nxt = (o_need_updat ? rsp_buf_ready_din : rsp_buf_ready_raw);
e603_subsys_gnrl_dfflrs  #(1) rsp_buf_ready_r_dfflrs    (rsp_buf_ready_r_ena, rsp_buf_ready_r_nxt, rsp_buf_ready_r,     clk, rst_n);// VPP_NO_REG_PARSE
  assign rsp_buf_ready = rsp_buf_ready_r;
  wire oo_outs_cnt_inc = o_icb_cmd_valid & o_icb_cmd_ready & o_clk_en 
                    ;
  wire oo_outs_cnt_dec = o_icb_rsp_valid & o_icb_rsp_ready & o_clk_en 
                    ;
  wire oo_outs_cnt_ena = oo_outs_cnt_inc ^ oo_outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] oo_outs_cnt_r;
  wire [OUTS_CNT_W-1:0] oo_outs_cnt_nxt = oo_outs_cnt_inc ? (oo_outs_cnt_r + 1'b1) : (oo_outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) oo_outs_cnt_dfflr (oo_outs_cnt_ena, oo_outs_cnt_nxt, oo_outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire oo_outs_cnt_eq0 = (oo_outs_cnt_r == {OUTS_CNT_W{1'b0}});
  assign oo_outs_cnt_max = (oo_outs_cnt_r == {OUTS_CNT_W{1'b1}});
  assign o_outs_cnt_max = (o_outs_cnt_r == {OUTS_CNT_W{1'b1}});
  if (RSP_STRICT_ORDER == 1) begin: rsp_strict_order_gen
      assign o_icb_rsp_valid_raw = (~oo_outs_cnt_eq0) & o_icb_rsp_valid;
      assign o_icb_rsp_ready     = (~oo_outs_cnt_eq0) & o_icb_rsp_ready_raw;
  end
  else begin: rsp_no_order_gen
      assign o_icb_rsp_valid_raw = o_icb_rsp_valid;
      assign o_icb_rsp_ready     = o_icb_rsp_ready_raw;
  end
  end
  endgenerate
endmodule
module e603_subsys_gnrl_ficb_async # (
    parameter RSP_STRICT_ORDER = 0,
  parameter PAYLOAD_NORST = 0,
  parameter RSP_ALWAYS_READY = 0,
  parameter OUTS_CNT_W = 1,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 4,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter AW = 32,
  parameter DW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  output             icb2icb_async_i_active,
  output             icb2icb_async_o_active,
  input              i_icb_cmd_sel  ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [DW-1:0]    i_icb_cmd_wdata,
  input  [DW/8-1:0]    i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [DW-1:0]    i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel  ,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [DW-1:0]    o_icb_cmd_wdata,
  output [DW/8-1:0]    o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input              i_clk,
  input              o_clk,
  input              i_rst_n,
  input              o_rst_n
  );
 wire i_icb_cmd_xlen_eq0 = (i_icb_cmd_xlen == 8'd0);
 wire i_icb_cmd_first = i_icb_cmd_beat[0] | i_icb_cmd_xlen_eq0;
 wire o_icb_cmd_xlen_eq0 = (o_icb_cmd_xlen == 8'd0);
 wire o_icb_cmd_first = o_icb_cmd_beat[0] | o_icb_cmd_xlen_eq0;
  wire i_icb_reset_flag_r;
e603_subsys_gnrl_dffrs #(1) reset_flag_dffrs (1'b0, i_icb_reset_flag_r, i_clk, i_rst_n);// VPP_NO_REG_PARSE
  localparam CMD_PACK_W = (1+AW+DW+DW/8+1+4+2+CMD_UW+8+2+2+1+3+0);
  wire [CMD_PACK_W-1:0] cmd_fifo_i_dat = {
                                 i_icb_cmd_read,
                                 i_icb_cmd_addr,
                                 i_icb_cmd_wdata,
                                 i_icb_cmd_wmask,
                                 i_icb_cmd_lock,
                                 i_icb_cmd_excl,
                                 i_icb_cmd_size,
                                 i_icb_cmd_beat,
                                 i_icb_cmd_xlen,
                                 i_icb_cmd_xburst,
                                 i_icb_cmd_modes,
                                 i_icb_cmd_dmode,
                                 i_icb_cmd_attri,
                                 i_icb_cmd_usr};
  wire [CMD_PACK_W-1:0] cmd_fifo_o_dat;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
    assign o_icb_cmd_size  = o_icb_cmd_size_pre ;
    assign o_icb_cmd_xlen  = o_icb_cmd_xlen_pre  ;
  assign {
                                 o_icb_cmd_read,
                                 o_icb_cmd_addr,
                                 o_icb_cmd_wdata,
                                 o_icb_cmd_wmask,
                                 o_icb_cmd_lock,
                                 o_icb_cmd_excl,
                                 o_icb_cmd_size_pre,
                                 o_icb_cmd_beat,
                                 o_icb_cmd_xlen_pre,
                                 o_icb_cmd_xburst,
                                 o_icb_cmd_modes,
                                 o_icb_cmd_dmode,
                                 o_icb_cmd_attri,
                                 o_icb_cmd_usr} = cmd_fifo_o_dat;
  wire cmd_fifo_i_valid;
  wire cmd_fifo_i_ready;
  wire outs_cnt_full;
  assign cmd_fifo_i_valid = (~i_icb_reset_flag_r) & (~outs_cnt_full) & i_icb_cmd_valid;
  assign i_icb_cmd_ready  = (~i_icb_reset_flag_r) & (~outs_cnt_full) & cmd_fifo_i_ready;
  wire o_icb_cmd_valid_pre;
  wire o_icb_cmd_ready_pre;
  wire i_cmd_cdc_active;
  wire o_cmd_cdc_active;
  wire i_rsp_cdc_active;
  wire o_rsp_cdc_active;
  generate
  if(ASYNC_FIFO == 0) begin: cdc_buf_cmd
  e603_subsys_gnrl_cdc_buf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DW     (CMD_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_buf_cmd(
    .i_clk    (i_clk),
    .i_rst_n  (i_rst_n),
    .i_vld    (cmd_fifo_i_valid),
    .i_rdy    (cmd_fifo_i_ready),
    .i_dat    (cmd_fifo_i_dat),
    .i_cdc_buf_active(i_cmd_cdc_active),
    .o_cdc_buf_active(o_cmd_cdc_active),
    .o_clk    (o_clk),
    .o_rst_n  (o_rst_n),
    .o_vld    (o_icb_cmd_valid_pre),
    .o_rdy    (o_icb_cmd_ready_pre),
    .o_dat    (cmd_fifo_o_dat )
  );
  end
  else begin: cdc_fifo_cmd
  e603_subsys_gnrl_cdc_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (CMD_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_cmd(
    .i_clk    (i_clk),
    .i_rst_n  (i_rst_n),
    .i_vld    (cmd_fifo_i_valid),
    .i_rdy    (cmd_fifo_i_ready),
    .i_dat    (cmd_fifo_i_dat),
    .i_cdc_fifo_active(i_cmd_cdc_active),
    .o_cdc_fifo_active(o_cmd_cdc_active),
    .o_clk    (o_clk),
    .o_rst_n  (o_rst_n),
    .o_vld    (o_icb_cmd_valid_pre),
    .o_rdy    (o_icb_cmd_ready_pre),
    .o_dat    (cmd_fifo_o_dat )
  );
  end
  endgenerate
  wire o_outs_cnt_max;
  wire rsp_buf_ready;
  generate
    if(RSP_ALWAYS_READY == 1) begin: gen_rsp_always_ready_1
      assign o_icb_cmd_valid     = rsp_buf_ready & o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = rsp_buf_ready & o_icb_cmd_ready;
    end
    else begin: gen_rsp_always_ready_0
      assign o_icb_cmd_valid     = o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = o_icb_cmd_ready;
    end
  endgenerate
  assign o_icb_cmd_sel = o_icb_cmd_valid_pre;
  localparam RSP_PACK_W = (2+DW+RSP_UW+0);
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata,
                                 o_icb_rsp_usr};
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 i_icb_rsp_err,
                                 i_icb_rsp_excl_ok,
                                 i_icb_rsp_rdata,
                                 i_icb_rsp_usr} = rsp_fifo_o_dat;
  wire o_icb_rsp_valid_raw;
  wire o_icb_rsp_ready_raw;
  generate
  if(ASYNC_FIFO == 0) begin: cdc_buf_rsp
  e603_subsys_gnrl_cdc_buf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DW     (RSP_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_buf_rsp(
    .i_clk    (o_clk),
    .i_rst_n  (o_rst_n),
    .i_vld   (o_icb_rsp_valid_raw),
    .i_rdy   (o_icb_rsp_ready_raw),
    .i_dat   (rsp_fifo_i_dat ),
    .i_cdc_buf_active(o_rsp_cdc_active),
    .o_cdc_buf_active(i_rsp_cdc_active),
    .o_clk    (i_clk),
    .o_rst_n  (i_rst_n),
    .o_vld  (i_icb_rsp_valid),
    .o_rdy  (i_icb_rsp_ready),
    .o_dat  (rsp_fifo_o_dat )
  );
  end
  else begin: cdc_fifo_rsp
  e603_subsys_gnrl_cdc_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP(ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (RSP_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_rsp(
    .i_clk    (o_clk),
    .i_rst_n  (o_rst_n),
    .i_vld   (o_icb_rsp_valid_raw),
    .i_rdy   (o_icb_rsp_ready_raw),
    .i_dat   (rsp_fifo_i_dat ),
    .i_cdc_fifo_active(o_rsp_cdc_active),
    .o_cdc_fifo_active(i_rsp_cdc_active),
    .o_clk    (i_clk),
    .o_rst_n  (i_rst_n),
    .o_vld  (i_icb_rsp_valid),
    .o_rdy  (i_icb_rsp_ready),
    .o_dat  (rsp_fifo_o_dat )
  );
  end
  endgenerate
  wire outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready
                    ;
  wire outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready
                    ;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, i_clk, i_rst_n);// VPP_NO_REG_PARSE
  assign outs_cnt_full = (outs_cnt_r == {OUTS_CNT_W{1'b1}});
  wire o_outs_cnt_inc = o_icb_cmd_valid & o_icb_cmd_ready 
                    ;
  wire o_outs_cnt_dec = o_icb_rsp_valid & o_icb_rsp_ready 
                    ;
  wire o_outs_cnt_ena = o_outs_cnt_inc ^ o_outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_r;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_nxt = o_outs_cnt_inc ? (o_outs_cnt_r + 1'b1) : (o_outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) o_outs_cnt_dfflr (o_outs_cnt_ena, o_outs_cnt_nxt, o_outs_cnt_r, o_clk, o_rst_n);// VPP_NO_REG_PARSE
  assign icb2icb_async_i_active = i_cmd_cdc_active | i_rsp_cdc_active | i_icb_cmd_valid | (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
  assign icb2icb_async_o_active = o_cmd_cdc_active | o_rsp_cdc_active | o_icb_cmd_valid_pre | (~(o_outs_cnt_r == {OUTS_CNT_W{1'b0}}));
  wire o_outs_cnt_eq0 = (o_outs_cnt_r == {OUTS_CNT_W{1'b0}});
  assign o_outs_cnt_max = (o_outs_cnt_r == {OUTS_CNT_W{1'b1}});
  generate
  if (RSP_STRICT_ORDER == 1) begin: rsp_strict_order_gen
      assign o_icb_rsp_valid_raw = (~o_outs_cnt_eq0) & o_icb_rsp_valid;
      assign o_icb_rsp_ready     = (~o_outs_cnt_eq0) & o_icb_rsp_ready_raw;
  end
  else begin: rsp_no_order_gen
      assign o_icb_rsp_valid_raw = o_icb_rsp_valid;
      assign o_icb_rsp_ready     = o_icb_rsp_ready_raw;
  end
  endgenerate
  assign rsp_buf_ready = (o_outs_cnt_r == {OUTS_CNT_W{1'b0}}) & o_icb_rsp_ready;
endmodule
module e603_subsys_gnrl_ficb_n2w # (
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 64
) (
  input              i_icb_cmd_sel ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
    wire cmd_y_lo_hi;
    wire rsp_y_lo_hi;
    wire rsp_y_lo_hi_real;
    wire rsp_y_merged;
    wire i_icb_rsp_hasked = i_icb_rsp_valid & i_icb_rsp_ready;
    assign rsp_y_lo_hi_real = rsp_y_lo_hi;
    wire i_icb_cmd_hasked = i_icb_cmd_valid & i_icb_cmd_ready;
    wire n2w_fifo_wen = o_icb_cmd_valid & o_icb_cmd_ready;
    wire n2w_fifo_ren = o_icb_rsp_valid & o_icb_rsp_ready;
    wire n2w_fifo_i_ready;
    wire n2w_fifo_i_valid = n2w_fifo_wen;
    wire n2w_fifo_full    = (~n2w_fifo_i_ready);
    wire n2w_fifo_o_valid ;
    wire n2w_fifo_o_ready = n2w_fifo_ren;
    wire n2w_fifo_empty   = (~n2w_fifo_o_valid);
    wire cmd_y_merged;
  generate
  if (ZEROCYC_RSP == 1) begin:gen_0cyc_rsp_1
      e603_subsys_gnrl_bypbuf #(
              .PAYLOAD_NORST(PAYLOAD_NORST),
              .DP  (FIFO_OUTS_NUM),
              .DW  (2)
      )  u_n2w_bypbuf(
          .i_vld(n2w_fifo_i_valid),
          .i_rdy(n2w_fifo_i_ready),
          .i_dat({cmd_y_lo_hi, cmd_y_merged} ),
          .o_dat({rsp_y_lo_hi, rsp_y_merged} ),
          .o_vld(n2w_fifo_o_valid),
          .o_rdy(n2w_fifo_o_ready),
          .fifo_o_vld(),
          .clk(clk),
          .rst_n(rst_n)
      );
  end
  else begin :gen_0cyc_rsp_0
      e603_subsys_gnrl_fifo # (
              .PAYLOAD_NORST(PAYLOAD_NORST),
        .CUT_READY (FIFO_CUT_READY),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
              .DW  (2)
      ) u_n2w_fifo (
        .i_vld(n2w_fifo_i_valid),
        .i_rdy(n2w_fifo_i_ready),
        .o_vld(n2w_fifo_o_valid),
        .o_rdy(n2w_fifo_o_ready),
          .i_dat({cmd_y_lo_hi, cmd_y_merged} ),
          .o_dat({rsp_y_lo_hi, rsp_y_merged} ),
        .clk  (clk),
        .rst_n(rst_n)
      );
  end
  endgenerate
  wire [AW-1:0]    i_icb_cmd_addr_algn;
  wire i_icb_cmd_size_full;
  wire i_icb_cmd_addr_lowr;
  generate
    if(X_W == 32) begin: gen_x_w_32
        assign cmd_y_lo_hi = i_icb_cmd_addr[2];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b10);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[2];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:3],3'b0};
    end
    if(X_W == 64) begin: gen_x_w_64
        assign cmd_y_lo_hi = i_icb_cmd_addr[3];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b11);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[3];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:4],4'b0};
    end
    if(X_W == 128) begin: gen_x_w_128
        assign cmd_y_lo_hi = i_icb_cmd_addr[4];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b100);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[4];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:5],5'b0};
    end
    if(X_W == 256) begin: gen_x_w_256
        assign cmd_y_lo_hi = i_icb_cmd_addr[5];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b101);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[5];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:6],6'b0};
    end
    if(X_W == 512) begin: gen_x_w_512
        assign cmd_y_lo_hi = i_icb_cmd_addr[6];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b110);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[6];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:7],7'b0};
    end
    if(X_W == 1024) begin: gen_x_w_1024
        assign cmd_y_lo_hi = i_icb_cmd_addr[7];
        assign i_icb_cmd_size_full = 1'b0;
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[7];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:8],8'b0};
    end
  endgenerate
  wire icb_2nd_flag_r;
  wire i_icb_cmd_fixed = (i_icb_cmd_xburst == 2'b00);
  wire i_icb_cmd_wrap = (i_icb_cmd_xburst == 2'b10);
  wire i_icb_cmd_wrap_xlen1 = i_icb_cmd_wrap & (~(| i_icb_cmd_xlen[7:1])) & i_icb_cmd_xlen[0];
  wire   i_icb_cmd_need_merg_pre =                    
                       (i_icb_cmd_xlen[0]) & 
                       i_icb_cmd_size_full &
                       ( i_icb_cmd_wrap_xlen1 ? 1'b1 : 
                                                i_icb_cmd_addr_lowr 
                       )
                       & (~i_icb_cmd_fixed)
                       ;
  wire   i_icb_cmd_need_merg = (~icb_2nd_flag_r) & i_icb_cmd_need_merg_pre;
  wire [Y_W-1:0]     o_icb_cmd_wdata_pre;
  wire [(Y_W/8-1):0] o_icb_cmd_wmask_pre;
  assign o_icb_cmd_wdata_pre = {i_icb_cmd_wdata,i_icb_cmd_wdata};
  assign o_icb_cmd_wmask_pre = cmd_y_lo_hi ?  {i_icb_cmd_wmask,  {X_W/8{1'b0}}} : {  {X_W/8{1'b0}},i_icb_cmd_wmask};
  wire i_icb_cmd_xlen_is1 = (i_icb_cmd_xlen == 8'd1);
  wire i_icb_cmd_xlen_is0 = (i_icb_cmd_xlen == 8'd0);
  wire i_cmd_xlen_cvt_incr = i_icb_cmd_xlen_is1 & i_icb_cmd_need_merg_pre;
  wire icb_2nd_cmd_valid_r;
  wire icb_2nd_cmd_read_r;
  wire i_icb_cmd_read_need_merg = 1'b0;
  assign cmd_y_merged = ( icb_2nd_cmd_valid_r 
                        )
                        ;
  wire o_icb_cmd_hasked  = o_icb_cmd_valid & o_icb_cmd_ready;
  wire n2w_icb_2nd_cmd_valid_set_raw = i_icb_cmd_need_merg & (~icb_2nd_cmd_valid_r); 
  wire n2w_icb_2nd_cmd_valid_set = n2w_icb_2nd_cmd_valid_set_raw & i_icb_cmd_hasked
             ;
  wire icb_2nd_cmd_valid_clr = o_icb_cmd_hasked & icb_2nd_cmd_valid_r;
  wire icb_2nd_cmd_valid_ena = n2w_icb_2nd_cmd_valid_set | icb_2nd_cmd_valid_clr;
  wire icb_2nd_cmd_valid_nxt = n2w_icb_2nd_cmd_valid_set;
e603_subsys_gnrl_dfflr #(1) icb_2nd_cmd_valid (icb_2nd_cmd_valid_ena, icb_2nd_cmd_valid_nxt, icb_2nd_cmd_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_2nd_flag_set = (~i_icb_cmd_xlen_is0) & i_icb_cmd_hasked & (~icb_2nd_flag_r) & (~i_icb_cmd_beat[1]);
  wire icb_2nd_flag_clr = i_icb_cmd_hasked & icb_2nd_flag_r;
  wire icb_2nd_flag_ena = icb_2nd_flag_set | icb_2nd_flag_clr;
  wire icb_2nd_flag_nxt = (~icb_2nd_flag_clr);
e603_subsys_gnrl_dfflr #(1) icb_2nd_flag (icb_2nd_flag_ena, icb_2nd_flag_nxt, icb_2nd_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire merg_buf_ena = n2w_icb_2nd_cmd_valid_set;
  wire [AW-1:0]    icb_2nd_cmd_addr_r;
  wire [X_W-1:0]   icb_2nd_cmd_wdata_r;
  wire [X_W/8-1:0] icb_2nd_cmd_wmask_r;
  wire             icb_2nd_cmd_beat0_r;
  wire i_icb_cmd_beat0 = i_icb_cmd_beat[0] & (~i_icb_cmd_xlen_is1);
e603_subsys_gnrl_dffl  #(AW)   icb_2nd_cmd_addr (merg_buf_ena, i_icb_cmd_addr_algn , icb_2nd_cmd_addr_r , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(X_W)  icb_2nd_cmd_wdata(merg_buf_ena, i_icb_cmd_wdata, icb_2nd_cmd_wdata_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(X_W/8)icb_2nd_cmd_wmask(merg_buf_ena, i_icb_cmd_wmask, icb_2nd_cmd_wmask_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)    icb_2nd_cmd_beat0(merg_buf_ena, i_icb_cmd_beat0 , icb_2nd_cmd_beat0_r , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)    icb_2nd_cmd_read (merg_buf_ena, i_icb_cmd_read  , icb_2nd_cmd_read_r  , clk, rst_n);// VPP_NO_REG_PARSE
  assign o_icb_cmd_sel   = (~n2w_fifo_full) & (i_icb_cmd_sel   | icb_2nd_cmd_valid_r);
  assign o_icb_cmd_valid = (~n2w_fifo_full) & (i_icb_cmd_need_merg ? (i_icb_cmd_valid & icb_2nd_cmd_valid_r) : i_icb_cmd_valid);
  assign i_icb_cmd_ready = (~n2w_fifo_full) & ((i_icb_cmd_need_merg & (~icb_2nd_cmd_valid_r)) ? 1'b1 : o_icb_cmd_ready);
  assign o_icb_cmd_addr  = 
            icb_2nd_cmd_valid_r ? icb_2nd_cmd_addr_r : i_icb_cmd_addr;
  assign o_icb_cmd_wdata = icb_2nd_cmd_valid_r ? (
                                 cmd_y_lo_hi ? {i_icb_cmd_wdata, icb_2nd_cmd_wdata_r} : {icb_2nd_cmd_wdata_r, i_icb_cmd_wdata}
                                 ) : o_icb_cmd_wdata_pre;
  assign o_icb_cmd_wmask = icb_2nd_cmd_valid_r ? (
                                 cmd_y_lo_hi ? {i_icb_cmd_wmask, icb_2nd_cmd_wmask_r} : {icb_2nd_cmd_wmask_r, i_icb_cmd_wmask}
                                 ) : o_icb_cmd_wmask_pre;
  wire             o_icb_cmd_read_pre;
  wire             o_icb_cmd_lock_pre;
  wire             o_icb_cmd_excl_pre;
  wire [1:0]       o_icb_cmd_modes_pre;
  wire             o_icb_cmd_dmode_pre;
  wire [1:0]       o_icb_cmd_xburst_pre;
  wire [2:0]       o_icb_cmd_attri_pre;
  assign o_icb_cmd_read_pre   = i_icb_cmd_read;
  assign o_icb_cmd_lock_pre   = i_icb_cmd_lock;
  assign o_icb_cmd_excl_pre   = i_icb_cmd_excl;
  assign o_icb_cmd_usr    = i_icb_cmd_usr;
  assign o_icb_cmd_xburst_pre = i_cmd_xlen_cvt_incr ? 2'b01 : i_icb_cmd_xburst;
  assign o_icb_cmd_modes_pre  = i_icb_cmd_modes ;
  assign o_icb_cmd_dmode_pre  = i_icb_cmd_dmode ;
  assign o_icb_cmd_attri_pre  = i_icb_cmd_attri ;
  assign o_icb_cmd_read   = o_icb_cmd_read_pre;
  assign o_icb_cmd_lock   = o_icb_cmd_lock_pre;
  assign o_icb_cmd_excl   = o_icb_cmd_excl_pre;
  assign o_icb_cmd_modes  = o_icb_cmd_modes_pre;
  assign o_icb_cmd_dmode  = o_icb_cmd_dmode_pre;
  assign o_icb_cmd_xburst = o_icb_cmd_xburst_pre;
  assign o_icb_cmd_attri  = o_icb_cmd_attri_pre;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
  wire [1:0] o_icb_cmd_beat_pre;
  assign o_icb_cmd_size = o_icb_cmd_size_pre;
  assign o_icb_cmd_xlen = o_icb_cmd_xlen_pre;
  assign o_icb_cmd_beat = o_icb_cmd_beat_pre;
  assign o_icb_cmd_beat_pre[0] = (icb_2nd_cmd_valid_r ? icb_2nd_cmd_beat0_r : i_icb_cmd_beat[0]) & (~i_cmd_xlen_cvt_incr);
  assign o_icb_cmd_beat_pre[1] = i_icb_cmd_beat[1] & (~(icb_2nd_cmd_valid_r & i_icb_cmd_xlen_is1));
  generate
  if (X_W == 32) begin:dw_64_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b011 : i_icb_cmd_size;
  end
  if (X_W == 64) begin:dw_128_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b100 : i_icb_cmd_size;
  end
  if (X_W == 128) begin:dw_256_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b101 : i_icb_cmd_size;
  end
  if (X_W == 256) begin:dw_512_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b110 : i_icb_cmd_size;
  end
  if (X_W == 512) begin:dw_1024_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b111 : i_icb_cmd_size;
  end
  if (X_W == 1024) begin:dw_2048_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b111 : i_icb_cmd_size;
  end
  endgenerate
    assign o_icb_cmd_xlen_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? {1'b0,i_icb_cmd_xlen[7:1]} : i_icb_cmd_xlen;
  wire icb_2nd_rsp_valid_r;
  wire icb_2nd_rsp_valid_set = (~icb_2nd_rsp_valid_r) & rsp_y_merged & i_icb_rsp_hasked;
  wire icb_2nd_rsp_valid_clr = icb_2nd_rsp_valid_r & i_icb_rsp_hasked;
  wire icb_2nd_rsp_valid_ena = icb_2nd_rsp_valid_set | icb_2nd_rsp_valid_clr;
  wire icb_2nd_rsp_valid_nxt = icb_2nd_rsp_valid_set;
e603_subsys_gnrl_dfflr #(1) icb_2nd_rsp_valid (icb_2nd_rsp_valid_ena, icb_2nd_rsp_valid_nxt, icb_2nd_rsp_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign o_icb_rsp_ready = (rsp_y_merged ? icb_2nd_rsp_valid_r : 1'b1) & i_icb_rsp_ready & n2w_fifo_o_valid;
  wire [X_W-1:0] i_icb_rsp_rdata_pre;
  wire [X_W-1:0] i_icb_rsp_rdata_merged;
  assign i_icb_rsp_rdata_pre    = rsp_y_lo_hi_real ? o_icb_rsp_rdata[Y_W-1:X_W] : o_icb_rsp_rdata[X_W-1:0] ;
  wire i_icb_rsp_rdata_merged_sel = (icb_2nd_rsp_valid_r ? rsp_y_lo_hi : (~rsp_y_lo_hi)); 
  assign i_icb_rsp_rdata_merged = i_icb_rsp_rdata_merged_sel 
                                     ? o_icb_rsp_rdata[Y_W-1:X_W] : o_icb_rsp_rdata[X_W-1:0] ;
  assign i_icb_rsp_rdata = rsp_y_merged ? i_icb_rsp_rdata_merged : i_icb_rsp_rdata_pre;
  assign i_icb_rsp_valid   = o_icb_rsp_valid & n2w_fifo_o_valid;  
  assign i_icb_rsp_err     = o_icb_rsp_err   ;
  assign i_icb_rsp_excl_ok = o_icb_rsp_excl_ok   ;
  assign i_icb_rsp_usr   = o_icb_rsp_usr   ;
endmodule
module e603_subsys_gnrl_ficb_nn2ww # (
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 128
) (
  input              i_icb_cmd_sel ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel  ,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W*2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W/4-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [7:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W*2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
  e603_subsys_gnrl_ficb_n2w # (
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W*2 )
  ) u_ficb_32to64 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel   ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_n2w # (
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W*2),
    .Y_W(Y_W )
  ) u_ficb_64to128 (
    .i_icb_cmd_sel       (dw_icb_cmd_sel  ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_nnn2www # (
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 128
) (
  input              i_icb_cmd_sel ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel  ,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W*2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W*2/8-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [7:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W*2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
  wire               dw2_icb_cmd_sel;
  wire               dw2_icb_cmd_valid;
  wire               dw2_icb_cmd_ready;
  wire               dw2_icb_cmd_read;
  wire [AW-1:0]      dw2_icb_cmd_addr;
  wire [X_W*4-1:0]      dw2_icb_cmd_wdata;
  wire [(X_W*4/8-1):0]  dw2_icb_cmd_wmask;
  wire               dw2_icb_cmd_lock;
  wire               dw2_icb_cmd_excl;
  wire [2:0]         dw2_icb_cmd_size;
  wire [1:0]         dw2_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw2_icb_cmd_usr;
  wire [7:0]         dw2_icb_cmd_xlen;
  wire [1:0]         dw2_icb_cmd_xburst;
  wire [1:0]         dw2_icb_cmd_modes;
  wire               dw2_icb_cmd_dmode;
  wire [2:0]         dw2_icb_cmd_attri;
  wire               dw2_icb_rsp_valid;
  wire               dw2_icb_rsp_ready;
  wire               dw2_icb_rsp_err;
  wire               dw2_icb_rsp_excl_ok;
  wire [X_W*4-1:0]      dw2_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw2_icb_rsp_usr;
  e603_subsys_gnrl_ficb_n2w # (
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W*2 )
  ) u_ficb_x_to_xm2 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel   ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_n2w # (
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W*2),
    .Y_W(X_W*4)
  ) u_ficb_xm2_to_xm4 (
    .i_icb_cmd_sel       (dw_icb_cmd_sel  ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .o_icb_cmd_sel       (dw2_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw2_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw2_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw2_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw2_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw2_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw2_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw2_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw2_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw2_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw2_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw2_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (dw2_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw2_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw2_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw2_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw2_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw2_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw2_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw2_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw2_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw2_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_n2w # (
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W*4),
    .Y_W(Y_W)
  ) u_ficb_xm4_to_y (
    .i_icb_cmd_sel       (dw2_icb_cmd_sel  ),
    .i_icb_cmd_valid     (dw2_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw2_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw2_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw2_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw2_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw2_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw2_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw2_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw2_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw2_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw2_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (dw2_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw2_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw2_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw2_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw2_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw2_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw2_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw2_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw2_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw2_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_w2n # (
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 64,
  parameter Y_W = 32
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  wire i_icb_rsp_err_pre;
  wire i_icb_rsp_excl_ok_pre;
  assign i_icb_rsp_err = i_icb_rsp_err_pre;
  assign i_icb_rsp_excl_ok = i_icb_rsp_excl_ok_pre;
  wire icb_cmd_size_dw;
  wire icb_cmd_addr_2 ;
  wire icb_cmd_size_dw_real = icb_cmd_size_dw;
generate
if (X_W == 64) begin:dw_64
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b11);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[2];
end
if (X_W == 128) begin:dw_128
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b100);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[3];
end
if (X_W == 256) begin:dw_256
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b101);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[4];
end
if (X_W == 512) begin:dw_512
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b110);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[5];
end
if (X_W == 1024) begin:dw_1024
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b111);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[6];
end
endgenerate
  wire o_icb_rsp_hasked  = o_icb_rsp_valid & o_icb_rsp_ready;
wire i_icb_cmd_fixed_cvt;
  wire w2n_fifo_wen = i_icb_cmd_valid & i_icb_cmd_ready;
  wire w2n_fifo_ren = i_icb_rsp_valid & i_icb_rsp_ready;
  wire w2n_fifo_i_valid = w2n_fifo_wen;
  wire w2n_fifo_i_ready;
  wire w2n_fifo_o_valid;
  wire w2n_fifo_o_match;
  wire w2n_has_ooo_id_buf;
  wire w2n_fifo_o_ready = w2n_fifo_ren;
  wire w2n_fifo_full;
    wire i_icb_cmd_xlen_is0 = (i_icb_cmd_xlen == {O_AXLEN_W{1'b0}});
    wire i_icb_xlen_overflow;
    wire icb_2nd_xlen_overflow;
    wire i_icb_cmd_xburst_fixed = (i_icb_cmd_xburst[1:0] == 2'b0);
    wire i_icb_cmd_xburst_fixed_xlen0     = (i_icb_cmd_xlen_is0 & i_icb_cmd_xburst_fixed);
    wire i_icb_cmd_xburst_fixed_n_xlen0 = ((~i_icb_cmd_xlen_is0) & i_icb_cmd_xburst_fixed);
    wire [1:0] i_icb_cmd_xburst_cvt = (i_icb_cmd_xburst_fixed_xlen0) ? 2'b01 : i_icb_cmd_xburst[1:0];
    assign i_icb_cmd_fixed_cvt = i_icb_cmd_xburst_fixed_n_xlen0 | i_icb_xlen_overflow; 
  wire icb_rsp_size_dw;
  wire icb_2nd_rsp_valid_r;
  wire o_icb_rsp_valid_dw = (icb_rsp_size_dw ? icb_2nd_rsp_valid_r : 1'b1);
  assign w2n_fifo_full = ~w2n_fifo_i_ready;
  wire w2n_fifo_empty = ~w2n_fifo_o_valid;
  wire icb_rsp_addr_2;
  wire icb_2nd_cmd_read_r;
  wire i_icb_cmd_last = i_icb_cmd_beat[1] | (i_icb_cmd_xlen == {O_AXLEN_W{1'b0}});
    wire icb_cmd_last = i_icb_cmd_last;
generate
if (ZEROCYC_RSP == 1) begin:gen_0cyc_rsp_1
    assign w2n_has_ooo_id_buf = 1'b0;
    assign w2n_fifo_o_match = 1'b0;
  e603_subsys_gnrl_bypbuf #(
    .PAYLOAD_NORST(PAYLOAD_NORST),
          .DP  (FIFO_OUTS_NUM),
          .DW  (2)
  )  u_rsp_w2n_bypbuf(
      .i_vld(w2n_fifo_i_valid),
      .i_rdy(w2n_fifo_i_ready),
      .i_dat({icb_cmd_size_dw_real,icb_cmd_addr_2}),
      .o_dat({icb_rsp_size_dw,icb_rsp_addr_2}),
      .o_vld(w2n_fifo_o_valid),
      .o_rdy(w2n_fifo_o_ready),
      .fifo_o_vld(),
      .clk(clk),
      .rst_n(rst_n)
  );
end
else begin :gen_0cyc_rsp_0
    if(SUPPORT_W2N_ID_OOO == 1) begin: id_ooo_is1
    assign w2n_has_ooo_id_buf = 1'b0;
    assign w2n_fifo_o_match = 1'b0;
      e603_subsys_gnrl_fifo #(
    .PAYLOAD_NORST(PAYLOAD_NORST),
          .CUT_READY (FIFO_CUT_READY),
          .MSKO      (0),
          .DW  (2),
          .DP  (FIFO_OUTS_NUM) 
      )  u_rsp_w2n_fifo(
          .i_vld(w2n_fifo_i_valid),
          .i_rdy(w2n_fifo_i_ready),
          .i_dat({icb_cmd_size_dw_real,icb_cmd_addr_2}),
          .o_dat({icb_rsp_size_dw,icb_rsp_addr_2}),
          .o_vld(w2n_fifo_o_valid),
          .o_rdy(w2n_fifo_o_ready),
          .clk(clk),
          .rst_n(rst_n)
      );
    end
    else begin: id_ooo_is0
    assign w2n_has_ooo_id_buf = 1'b0;
    assign w2n_fifo_o_match = 1'b0;
      e603_subsys_gnrl_fifo #(
    .PAYLOAD_NORST(PAYLOAD_NORST),
          .CUT_READY (FIFO_CUT_READY),
          .MSKO      (0),
          .DP  (FIFO_OUTS_NUM),
          .DW  (2)
      )  u_rsp_w2n_fifo(
          .i_vld(w2n_fifo_i_valid),
          .i_rdy(w2n_fifo_i_ready),
          .i_dat({icb_cmd_size_dw_real,icb_cmd_addr_2}),
          .o_dat({icb_rsp_size_dw,icb_rsp_addr_2}),
          .o_vld(w2n_fifo_o_valid),
          .o_rdy(w2n_fifo_o_ready),
          .clk(clk),
          .rst_n(rst_n)
      );
    end
end
endgenerate
  wire             icb_2nd_cmd_valid_r;
  wire             icb_2nd_cmd_valid_ena;
  wire             icb_2nd_cmd_valid_nxt;
  wire             icb_2nd_cmd_valid_set;
  wire             icb_2nd_cmd_valid_clr;
  wire             i_icb_cmd_ready_addi_cond;
  wire o_icb_cmd_hasked  = o_icb_cmd_valid & o_icb_cmd_ready;
    wire i_icb_cvt_single;
    wire icb_2nd_cmd_valid_set_raw     = icb_cmd_size_dw      & o_icb_cmd_hasked & (~icb_2nd_cmd_valid_r);
    assign icb_2nd_cmd_valid_set     = icb_2nd_cmd_valid_set_raw;
    wire icb_2nd_cmd_set = icb_2nd_cmd_valid_set;
    assign icb_2nd_cmd_valid_clr     = icb_2nd_cmd_valid_r  & o_icb_cmd_hasked;
    wire icb_2nd_cmd_valid_real;
    assign icb_2nd_cmd_valid_real = icb_2nd_cmd_valid_r;
    assign i_icb_cmd_ready_addi_cond = !icb_2nd_cmd_valid_real;
    assign i_icb_cmd_ready = (~w2n_fifo_full) & i_icb_cmd_ready_addi_cond & o_icb_cmd_ready;
    wire             icb_2nd_cmd_excl_r;
    wire             icb_2nd_cmd_lock_r;
    wire [AW-1:0]    icb_2nd_cmd_addr_r;
    wire [Y_W-1:0]   icb_2nd_cmd_wdata_r;
    wire [Y_W/8-1:0] icb_2nd_cmd_wmask_r;
    wire [CMD_UW-1:0] icb_2nd_cmd_usr_r;
    wire [1:0] icb_2nd_cmd_beat_r;
    wire [O_AXLEN_W-1:0] icb_2nd_cmd_xlen_r  ;
    wire [1:0] icb_2nd_cmd_xburst_r;
    wire [1:0] icb_2nd_cmd_modes_r ;
    wire icb_2nd_load_ena = icb_2nd_cmd_set;
    wire       icb_2nd_cmd_dmode_r ;
    wire [2:0] icb_2nd_cmd_attri_r ;
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_lock   (icb_2nd_load_ena, i_icb_cmd_lock, icb_2nd_cmd_lock_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_excl   (icb_2nd_load_ena, i_icb_cmd_excl, icb_2nd_cmd_excl_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_read   (icb_2nd_load_ena, i_icb_cmd_read, icb_2nd_cmd_read_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(AW)  icb_2nd_cmd_addr   (icb_2nd_cmd_set, i_icb_cmd_addr[AW-1:0], icb_2nd_cmd_addr_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(Y_W)   icb_2nd_cmd_wdata  (icb_2nd_load_ena, i_icb_cmd_wdata[X_W-1:Y_W], icb_2nd_cmd_wdata_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(Y_W/8) icb_2nd_cmd_wmask  (icb_2nd_load_ena, i_icb_cmd_wmask[X_W/8-1:Y_W/8], icb_2nd_cmd_wmask_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(CMD_UW)icb_2nd_cmd_usr    (icb_2nd_load_ena, i_icb_cmd_usr, icb_2nd_cmd_usr_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2)     icb_2nd_cmd_beat   (icb_2nd_load_ena, i_icb_cmd_beat, icb_2nd_cmd_beat_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(O_AXLEN_W)     icb_2nd_cmd_xlen   (icb_2nd_load_ena, i_icb_cmd_xlen  , icb_2nd_cmd_xlen_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2)     icb_2nd_cmd_xburst (icb_2nd_load_ena, i_icb_cmd_xburst_cvt, icb_2nd_cmd_xburst_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2)     icb_2nd_cmd_modes  (icb_2nd_load_ena, i_icb_cmd_modes , icb_2nd_cmd_modes_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_dmode  (icb_2nd_load_ena, i_icb_cmd_dmode , icb_2nd_cmd_dmode_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(3)     icb_2nd_cmd_attri  (icb_2nd_load_ena, i_icb_cmd_attri , icb_2nd_cmd_attri_r, clk, rst_n);// VPP_NO_REG_PARSE
    assign o_icb_cmd_sel   = (~w2n_fifo_full) & i_icb_cmd_sel   || icb_2nd_cmd_valid_real;
    assign o_icb_cmd_valid = (~w2n_fifo_full) & i_icb_cmd_valid || icb_2nd_cmd_valid_real;
  wire [2:0] o_icb_cmd_size_pre;
  wire [O_AXLEN_W-1:0] o_icb_cmd_xlen_pre;
  wire [1:0] o_icb_cmd_beat_pre;
  wire [AW-1:0] o_icb_cmd_addr_pre;
  assign o_icb_cmd_size = o_icb_cmd_size_pre;
  assign o_icb_cmd_xlen = o_icb_cmd_xlen_pre;
  assign o_icb_cmd_beat = o_icb_cmd_beat_pre;
  assign o_icb_cmd_addr = o_icb_cmd_addr_pre;
  wire             o_icb_cmd_read_pre;
  wire             o_icb_cmd_lock_pre;
  wire             o_icb_cmd_excl_pre;
  wire [1:0]       o_icb_cmd_modes_pre;
  wire             o_icb_cmd_dmode_pre;
  wire [1:0]       o_icb_cmd_xburst_pre;
  wire [2:0]       o_icb_cmd_attri_pre;
  assign o_icb_cmd_read   = o_icb_cmd_read_pre;
  assign o_icb_cmd_lock   = o_icb_cmd_lock_pre;
  assign o_icb_cmd_excl   = o_icb_cmd_excl_pre;
  assign o_icb_cmd_modes  = o_icb_cmd_modes_pre ;
  assign o_icb_cmd_dmode  = o_icb_cmd_dmode_pre ;
  assign o_icb_cmd_attri  = o_icb_cmd_attri_pre ;
  assign o_icb_cmd_xburst = o_icb_cmd_xburst_pre ;
    assign o_icb_cmd_addr_pre = icb_2nd_cmd_valid_r ? (
                                                    (X_W == 64) ? {icb_2nd_cmd_addr_r[AW-1:3],3'b100} :
                                                    (X_W == 256) ? {icb_2nd_cmd_addr_r[AW-1:5],5'b10000} :
                                                    (X_W == 512) ? {icb_2nd_cmd_addr_r[AW-1:6],6'b100000} :
                                                    (X_W == 1024) ? {icb_2nd_cmd_addr_r[AW-1:7],7'b1000000} :
                                                                  {icb_2nd_cmd_addr_r[AW-1:4],4'b1000}
                                                    ) :
                             icb_cmd_size_dw    ? (
                                                    (X_W == 64) ? {i_icb_cmd_addr[AW-1:3],3'b0} :
                                                    (X_W == 256) ? {i_icb_cmd_addr[AW-1:5],5'b0} :
                                                    (X_W == 512) ? {i_icb_cmd_addr[AW-1:6],6'b0} :
                                                    (X_W == 1024) ? {i_icb_cmd_addr[AW-1:7],7'b0} :
                                                                  {i_icb_cmd_addr[AW-1:4],4'b0}
                                                    )
                                                :  i_icb_cmd_addr;
    assign o_icb_cmd_read_pre = icb_2nd_cmd_valid_real ? icb_2nd_cmd_read_r
                                                : i_icb_cmd_read;
    assign o_icb_cmd_lock_pre = icb_2nd_cmd_valid_real ? icb_2nd_cmd_lock_r
                                                : i_icb_cmd_lock;
    assign o_icb_cmd_excl_pre = icb_2nd_cmd_valid_real ? icb_2nd_cmd_excl_r
                                                : i_icb_cmd_excl;
    assign o_icb_cmd_wdata = icb_2nd_cmd_valid_real ? icb_2nd_cmd_wdata_r :
                             icb_cmd_size_dw     ? i_icb_cmd_wdata[Y_W-1:0] :
                             icb_cmd_addr_2      ? i_icb_cmd_wdata[X_W-1:Y_W] :
                                                   i_icb_cmd_wdata[Y_W-1:0];
    assign o_icb_cmd_wmask = icb_2nd_cmd_valid_real ? icb_2nd_cmd_wmask_r :
                             icb_cmd_size_dw     ? i_icb_cmd_wmask[(Y_W/8-1):0] :
                             icb_cmd_addr_2      ? i_icb_cmd_wmask[(X_W/8-1):(Y_W/8)] :
                                                   i_icb_cmd_wmask[(Y_W/8-1):0];
    assign o_icb_cmd_usr  = icb_2nd_cmd_valid_real ? icb_2nd_cmd_usr_r : i_icb_cmd_usr;
  generate
    if(O_AXLEN_EXTEND == 1) begin: xlen_extend_1_gen
        assign i_icb_xlen_overflow   = 1'b0;
        assign icb_2nd_xlen_overflow = 1'b0;
    end
    else begin: xlen_extend_0_gen
        assign i_icb_xlen_overflow = 
                    (icb_cmd_size_dw & (i_icb_cmd_xburst == 2'b10)) ? i_icb_cmd_xlen[3] : 
                    (icb_cmd_size_dw & (i_icb_cmd_xburst == 2'b01)) ? i_icb_cmd_xlen[7] : 1'b0 ;
        assign icb_2nd_xlen_overflow= (
                   (icb_2nd_cmd_xburst_r == 2'b10) ? icb_2nd_cmd_xlen_r[3] :
                   (icb_2nd_cmd_xburst_r == 2'b01) ? icb_2nd_cmd_xlen_r[7] : 1'b0) ;
    end
  endgenerate
    wire icb_2nd_cvt_single = (icb_2nd_cmd_xburst_r == 2'b0) | icb_2nd_xlen_overflow;
    assign i_icb_cvt_single   = i_icb_cmd_fixed_cvt;
    wire icb_2nd_cmd_xlen_is0 = (icb_2nd_cmd_xlen_r == {O_AXLEN_W{1'd0}});
    assign o_icb_cmd_beat_pre[0] = icb_2nd_cmd_valid_r ? (1'b0                                                                    ) : ((~i_icb_cvt_single) & (i_icb_cmd_beat[0] | (icb_cmd_size_dw & i_icb_cmd_xlen_is0)));
    assign o_icb_cmd_beat_pre[1] = icb_2nd_cmd_valid_r ? ((~icb_2nd_cvt_single) & (icb_2nd_cmd_beat_r[1] | (icb_2nd_cmd_xlen_is0))) : ((~i_icb_cvt_single) & (icb_cmd_size_dw ? 1'b0 : i_icb_cmd_beat[1]));
    wire [O_AXLEN_W-1:0] o_icb_cmd_xlen_raw;
    generate
    if (X_W == 64) begin:dw_64_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b10 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 128) begin:dw_128_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b11 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 256) begin:dw_256_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b100: i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 512) begin:dw_512_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b101 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 1024) begin:dw_1024_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b110 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    endgenerate
    assign o_icb_cmd_xlen_pre = o_icb_cmd_xlen_raw;
    assign o_icb_cmd_xburst_pre  = icb_2nd_cmd_valid_real ? (icb_2nd_cvt_single ? 2'b01 : icb_2nd_cmd_xburst_r)
                                                   : (i_icb_cvt_single ? 2'b01 : i_icb_cmd_xburst_cvt);
    assign o_icb_cmd_modes_pre   = icb_2nd_cmd_valid_real ? icb_2nd_cmd_modes_r  : i_icb_cmd_modes ;
    assign o_icb_cmd_dmode_pre   = icb_2nd_cmd_valid_real ? icb_2nd_cmd_dmode_r  : i_icb_cmd_dmode ;
    assign o_icb_cmd_attri_pre   = icb_2nd_cmd_valid_real ? icb_2nd_cmd_attri_r  : i_icb_cmd_attri ;
  assign icb_2nd_cmd_valid_ena = icb_2nd_cmd_valid_set | icb_2nd_cmd_valid_clr;
  assign icb_2nd_cmd_valid_nxt = icb_2nd_cmd_valid_set & (~icb_2nd_cmd_valid_clr);
e603_subsys_gnrl_dfflr #(1)     icb_2nd_cmd_valid  (icb_2nd_cmd_valid_ena, icb_2nd_cmd_valid_nxt, icb_2nd_cmd_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire i_icb_rsp_hasked  = i_icb_rsp_valid & i_icb_rsp_ready;
  wire icb_2nd_rsp_valid_set = icb_rsp_size_dw & o_icb_rsp_hasked & (~icb_2nd_rsp_valid_r);
  wire icb_2nd_rsp_valid_clr = icb_rsp_size_dw & o_icb_rsp_hasked & icb_2nd_rsp_valid_r;
  wire icb_2nd_rsp_valid_ena = icb_2nd_rsp_valid_set | icb_2nd_rsp_valid_clr;
  wire icb_2nd_rsp_valid_nxt = icb_2nd_rsp_valid_set & (~icb_2nd_rsp_valid_clr);
e603_subsys_gnrl_dfflr #(1) icb_2nd_rsp_valid_dfflr(icb_2nd_rsp_valid_ena, icb_2nd_rsp_valid_nxt, icb_2nd_rsp_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_ena = icb_rsp_size_dw &  o_icb_rsp_hasked & (~icb_2nd_rsp_valid_r);
  wire [Y_W-1:0] icb_rsp_leftover_rdata_nxt = o_icb_rsp_rdata[Y_W-1:0];
  wire [Y_W-1:0] icb_rsp_leftover_rdata_r;
e603_subsys_gnrl_dffl  #(Y_W) icb_rsp_leftover_rdata_dffl (icb_rsp_leftover_ena, icb_rsp_leftover_rdata_nxt, icb_rsp_leftover_rdata_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_err_nxt = o_icb_rsp_err;
  wire icb_rsp_leftover_err_r;
e603_subsys_gnrl_dffl  #(1) icb_rsp_leftover_err_dffl (icb_rsp_leftover_ena, icb_rsp_leftover_err_nxt, icb_rsp_leftover_err_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_excl_ok_nxt = o_icb_rsp_excl_ok;
  wire icb_rsp_leftover_excl_ok_r;
e603_subsys_gnrl_dffl  #(1) icb_rsp_leftover_excl_ok_dffl                   (icb_rsp_leftover_ena, icb_rsp_leftover_excl_ok_nxt, icb_rsp_leftover_excl_ok_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_vld = icb_2nd_rsp_valid_r;
  wire i_icb_rsp_valid_cond = (icb_rsp_size_dw ? icb_2nd_rsp_valid_r : 1'b1)
                            ;
  wire o_icb_rsp_ready_byp = (icb_rsp_size_dw & (~icb_2nd_rsp_valid_r))
                             ;
  wire w2n_fifo_o_valid_real = w2n_has_ooo_id_buf ? w2n_fifo_o_match : w2n_fifo_o_valid;
  assign i_icb_rsp_valid =  i_icb_rsp_valid_cond & o_icb_rsp_valid & w2n_fifo_o_valid_real;
  assign i_icb_rsp_rdata = icb_rsp_leftover_vld ? {o_icb_rsp_rdata, icb_rsp_leftover_rdata_r} :
                           icb_rsp_addr_2       ? {o_icb_rsp_rdata, {Y_W{1'b0}}}              :
                                                  {{Y_W{1'b0}}, o_icb_rsp_rdata}
                                                ;
  assign o_icb_rsp_ready = (o_icb_rsp_ready_byp ? 1'b1 : i_icb_rsp_ready) & w2n_fifo_o_valid_real;
  assign i_icb_rsp_err_pre   = icb_rsp_leftover_vld ? (|{icb_rsp_leftover_err_r, o_icb_rsp_err
                                                          }) : 
                                                             (|{
                                                              o_icb_rsp_err
                                                              });
  assign i_icb_rsp_excl_ok_pre = icb_rsp_leftover_vld ? |{icb_rsp_leftover_excl_ok_r, o_icb_rsp_excl_ok} : o_icb_rsp_excl_ok;
  assign i_icb_rsp_usr   = o_icb_rsp_usr;
endmodule
module e603_subsys_gnrl_ficb_ww2nn # (
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 0,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 128,
  parameter Y_W = 32
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W/2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W/16-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [O_AXLEN_W-1:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W/2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
  e603_subsys_gnrl_ficb_w2n # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W/2 )
  ) u_ficb_x2x_div2 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_w2n # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W/2),
    .Y_W(Y_W )
  ) u_ficb_x_div2_to_y (
    .i_icb_cmd_sel       (dw_icb_cmd_sel    ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_www2nnn # (
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 0,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 256,
  parameter Y_W = 32
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W/2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W/16-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [O_AXLEN_W-1:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W/2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
 wire                dw2_icb_cmd_sel;
  wire               dw2_icb_cmd_valid;
  wire               dw2_icb_cmd_ready;
  wire               dw2_icb_cmd_read;
  wire [AW-1:0]      dw2_icb_cmd_addr;
  wire [X_W/4-1:0]   dw2_icb_cmd_wdata;
  wire [(X_W/32-1):0]dw2_icb_cmd_wmask;
  wire               dw2_icb_cmd_lock;
  wire               dw2_icb_cmd_excl;
  wire [2:0]         dw2_icb_cmd_size;
  wire [1:0]         dw2_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw2_icb_cmd_usr;
  wire [O_AXLEN_W-1:0]         dw2_icb_cmd_xlen;
  wire [1:0]         dw2_icb_cmd_xburst;
  wire [1:0]         dw2_icb_cmd_modes;
  wire               dw2_icb_cmd_dmode;
  wire [2:0]         dw2_icb_cmd_attri;
  wire               dw2_icb_rsp_valid;
  wire               dw2_icb_rsp_ready;
  wire               dw2_icb_rsp_err;
  wire               dw2_icb_rsp_excl_ok;
  wire [X_W/4-1:0]   dw2_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw2_icb_rsp_usr;
  e603_subsys_gnrl_ficb_w2n # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W/2 )
  ) u_ficb_x2x_div2 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_w2n # (
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W/2),
    .Y_W(X_W/4)
  ) u_ficb_x_div2_to_x_div4 (
    .i_icb_cmd_sel       (dw_icb_cmd_sel    ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .o_icb_cmd_sel       (dw2_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw2_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw2_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw2_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw2_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw2_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw2_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw2_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw2_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw2_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw2_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw2_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (dw2_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw2_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw2_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw2_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw2_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw2_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw2_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw2_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw2_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw2_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_w2n # (
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W/4),
    .Y_W(Y_W)
  ) u_ficb_x_div4_to_y (
    .i_icb_cmd_sel       (dw2_icb_cmd_sel    ),
    .i_icb_cmd_valid     (dw2_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw2_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw2_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw2_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw2_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw2_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw2_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw2_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw2_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw2_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw2_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (dw2_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw2_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw2_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw2_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw2_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw2_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw2_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw2_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw2_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw2_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_wconv # (
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 0,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter RSP_CHECK_CMD_OUTS = 0,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 64
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  generate
    if(X_W == Y_W) begin: x_is_y_gen
    wire rspid_fifo_i_ready;
    wire rspid_fifo_o_valid;
        if(RSP_CHECK_CMD_OUTS == 1) begin: rsp_fifo_gen
    wire rspid_fifo_i_push = o_icb_cmd_valid & o_icb_cmd_ready
                           ;
    wire rspid_fifo_o_pop  = o_icb_rsp_valid & o_icb_rsp_ready
                           ;
    e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT(1'b1),
        .CUT_READY (FIFO_CUT_READY),
        .DP  (FIFO_OUTS_NUM+1),
        .DW  (1)
      ) u_e603_subsys_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_push ),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(1'b0 ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_pop),
        .o_dat(),
        .clk  (clk),
        .rst_n(rst_n)
      );
        end
        else begin : no_rsp_fifo_gen
    assign rspid_fifo_i_ready = 1'b1;
    assign rspid_fifo_o_valid = 1'b1;
        end
        assign o_icb_cmd_sel   = i_icb_cmd_sel;
        assign i_icb_cmd_ready = rspid_fifo_i_ready & o_icb_cmd_ready;
        assign o_icb_cmd_valid = rspid_fifo_i_ready & i_icb_cmd_valid;
        assign o_icb_cmd_read  = i_icb_cmd_read ;
        assign o_icb_cmd_addr  = i_icb_cmd_addr ;
        assign o_icb_cmd_wdata = i_icb_cmd_wdata;
        assign o_icb_cmd_wmask = i_icb_cmd_wmask;
        assign o_icb_cmd_beat  = i_icb_cmd_beat ;
        assign o_icb_cmd_lock  = i_icb_cmd_lock ;
        assign o_icb_cmd_excl  = i_icb_cmd_excl ;
        assign o_icb_cmd_size  = i_icb_cmd_size ;
        assign o_icb_cmd_usr   = i_icb_cmd_usr  ;
        assign o_icb_cmd_xlen  = i_icb_cmd_xlen  ;
        assign o_icb_cmd_xburst= i_icb_cmd_xburst;
        assign o_icb_cmd_modes = i_icb_cmd_modes ;
        assign o_icb_cmd_dmode = i_icb_cmd_dmode ;
        assign o_icb_cmd_attri = i_icb_cmd_attri ;
        assign o_icb_rsp_ready     = rspid_fifo_o_valid & i_icb_rsp_ready;
        assign i_icb_rsp_valid     = rspid_fifo_o_valid & o_icb_rsp_valid;
        assign i_icb_rsp_err       = o_icb_rsp_err  ;
        assign i_icb_rsp_excl_ok   = o_icb_rsp_excl_ok  ;
        assign i_icb_rsp_rdata     = o_icb_rsp_rdata;
        assign i_icb_rsp_usr       = o_icb_rsp_usr;
    end
    if(    ((Y_W ==  64) && (X_W ==  32)) 
        || ((Y_W == 128) && (X_W ==  64))
        || ((Y_W == 256) && (X_W == 128))
        || ((Y_W == 512) && (X_W == 256))
        || ((Y_W == 1024) && (X_W == 512))
        || ((Y_W == 2048) && (X_W == 1024))
        ) begin:n2w_gen
  e603_subsys_gnrl_ficb_n2w # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_n2w (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((Y_W == 128) && (X_W == 32))
      || ((Y_W == 256) && (X_W == 64))
      || ((Y_W == 512) && (X_W == 128))
      || ((Y_W == 1024) && (X_W == 256))
      || ((Y_W == 2048) && (X_W == 512))
        ) begin:nn2ww_gen
  e603_subsys_gnrl_ficb_nn2ww # (
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_nn2ww (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((Y_W == 256) && (X_W == 32))
      || ((Y_W == 512) && (X_W == 64))
      || ((Y_W == 1024) && (X_W == 128))
      || ((Y_W == 2048) && (X_W == 256))
        ) begin:nnn2www_gen
  e603_subsys_gnrl_ficb_nnn2www # (
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_nnn2www (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(    ((X_W ==  64) && (Y_W ==  32)) 
        || ((X_W == 128) && (Y_W ==  64))
        || ((X_W == 256) && (Y_W == 128))
        || ((X_W == 512) && (Y_W == 256))
        || ((X_W == 1024) && (Y_W == 512))
        ) begin:w2n_gen
  e603_subsys_gnrl_ficb_w2n # (
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_w2n (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((X_W == 128) && (Y_W == 32))
      || ((X_W == 256) && (Y_W == 64))
      || ((X_W == 512) && (Y_W == 128))
      || ((X_W == 1024) && (Y_W == 256))
        ) begin:ww2nn
  e603_subsys_gnrl_ficb_ww2nn # (
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_ww2nn (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((X_W == 256) && (Y_W == 32))
      || ((X_W == 512) && (Y_W == 64))
      || ((X_W == 1024) && (Y_W == 128))
        ) begin:www2nnn
  e603_subsys_gnrl_ficb_www2nnn # (
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_www2nnn (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
  endgenerate
endmodule
module e603_subsys_gnrl_ficb_splt
 # (
  parameter AW = 32,
  parameter DW = 64,
  parameter USE_ALL_READY = 0,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter SPLT_NUM = 4,
  parameter SPLT_PTR_1HOT = 1,
  parameter PAYLOAD_NORST = 0,
  parameter SPLT_PTR_W = 4,
  parameter FIFO_REG_OUT = 0,
  parameter ALLOW_DIFF = 1,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  input  [SPLT_NUM-1:0] i_icb_splt_indic,
  output splt_active,
  input  clk_en,
  input  i_icb_cmd_sel,
  input  i_icb_cmd_valid,
  output i_icb_cmd_ready,
  input             i_icb_cmd_read,
  input  [AW-1:0]   i_icb_cmd_addr,
  input  [DW-1:0]   i_icb_cmd_wdata,
  input  [DW/8-1:0]   i_icb_cmd_wmask,
  input  [1:0]      i_icb_cmd_beat,
  input             i_icb_cmd_lock,
  input             i_icb_cmd_excl,
  input  [2:0]      i_icb_cmd_size,
  input  [CMD_UW-1:0]i_icb_cmd_usr,
  input [7:0]       i_icb_cmd_xlen,
  input [1:0]       i_icb_cmd_xburst,
  input [1:0]       i_icb_cmd_modes,
  input             i_icb_cmd_dmode,
  input [2:0]       i_icb_cmd_attri,
  output i_icb_rsp_valid,
  input  i_icb_rsp_ready,
  output i_icb_rsp_err,
  output i_icb_rsp_excl_ok,
  output [DW-1:0] i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  input  [SPLT_NUM*1-1:0]    o_bus_icb_cmd_ready,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_valid,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_sel,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_read,
  output [SPLT_NUM*AW-1:0]   o_bus_icb_cmd_addr,
  output [SPLT_NUM*DW-1:0]   o_bus_icb_cmd_wdata,
  output [SPLT_NUM*DW/8-1:0]   o_bus_icb_cmd_wmask,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_beat,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_lock,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_excl,
  output [SPLT_NUM*3-1:0]    o_bus_icb_cmd_size,
  output [SPLT_NUM*CMD_UW-1:0]o_bus_icb_cmd_usr,
  output [SPLT_NUM*8-1:0]    o_bus_icb_cmd_xlen,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_xburst,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_modes,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_dmode,
  output [SPLT_NUM*3-1:0]    o_bus_icb_cmd_attri,
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_valid,
  output [SPLT_NUM*1-1:0]  o_bus_icb_rsp_ready,
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_err,
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_excl_ok,
  input  [SPLT_NUM*DW-1:0] o_bus_icb_rsp_rdata,
  input  [SPLT_NUM*RSP_UW-1:0] o_bus_icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  wire [SPLT_NUM-1:0] i_icb_splt_indic_real;
    wire i_icb_cmd_hsked = i_icb_cmd_valid & i_icb_cmd_ready;
    assign i_icb_splt_indic_real = i_icb_splt_indic;
  localparam SPLT_FIFO_DW = SPLT_PTR_W 
                       ;
  wire rspid_fifo_empty;
generate 
  if(SPLT_NUM == 1) begin:gen_splt_num_eq_1
    assign i_icb_cmd_ready     = o_bus_icb_cmd_ready;
    assign o_bus_icb_cmd_sel   = i_icb_cmd_sel;
    assign o_bus_icb_cmd_valid = i_icb_cmd_valid;
    assign o_bus_icb_cmd_read  = i_icb_cmd_read ;
    assign o_bus_icb_cmd_addr  = i_icb_cmd_addr ;
    assign o_bus_icb_cmd_wdata = i_icb_cmd_wdata;
    assign o_bus_icb_cmd_wmask = i_icb_cmd_wmask;
    assign o_bus_icb_cmd_beat  = i_icb_cmd_beat ;
    assign o_bus_icb_cmd_lock  = i_icb_cmd_lock ;
    assign o_bus_icb_cmd_excl  = i_icb_cmd_excl ;
    assign o_bus_icb_cmd_size  = i_icb_cmd_size ;
    assign o_bus_icb_cmd_usr   = i_icb_cmd_usr  ;
    assign o_bus_icb_cmd_xlen  = i_icb_cmd_xlen  ;
    assign o_bus_icb_cmd_xburst= i_icb_cmd_xburst;
    assign o_bus_icb_cmd_modes = i_icb_cmd_modes ;
    assign o_bus_icb_cmd_dmode = i_icb_cmd_dmode ;
    assign o_bus_icb_cmd_attri = i_icb_cmd_attri ;
    assign rspid_fifo_empty    = 1'b1;
    assign o_bus_icb_rsp_ready = i_icb_rsp_ready;
    assign i_icb_rsp_valid     = o_bus_icb_rsp_valid;
    assign i_icb_rsp_err       = o_bus_icb_rsp_err  ;
    assign i_icb_rsp_excl_ok   = o_bus_icb_rsp_excl_ok  ;
    assign i_icb_rsp_rdata     = o_bus_icb_rsp_rdata;
    assign i_icb_rsp_usr       = o_bus_icb_rsp_usr;
  end
  else begin:gen_splt_num_gt_1
    genvar i;
    genvar ii;
    integer j;
    wire [SPLT_NUM-1:0] o_icb_cmd_sel;
    wire [SPLT_NUM-1:0] o_icb_cmd_valid;
    wire [SPLT_NUM-1:0] o_icb_cmd_ready;
    wire            o_icb_cmd_read [SPLT_NUM-1:0];
    wire [AW-1:0]   o_icb_cmd_addr [SPLT_NUM-1:0];
    wire [DW-1:0]   o_icb_cmd_wdata[SPLT_NUM-1:0];
    wire [DW/8-1:0]   o_icb_cmd_wmask[SPLT_NUM-1:0];
    wire [1:0]      o_icb_cmd_beat [SPLT_NUM-1:0];
    wire            o_icb_cmd_lock [SPLT_NUM-1:0];
    wire            o_icb_cmd_excl [SPLT_NUM-1:0];
    wire [2:0]      o_icb_cmd_size [SPLT_NUM-1:0];
    wire [CMD_UW-1:0]o_icb_cmd_usr  [SPLT_NUM-1:0];
    wire [7:0]      o_icb_cmd_xlen  [SPLT_NUM-1:0];
    wire [1:0]      o_icb_cmd_xburst[SPLT_NUM-1:0];
    wire [1:0]      o_icb_cmd_modes [SPLT_NUM-1:0];
    wire            o_icb_cmd_dmode [SPLT_NUM-1:0];
    wire [2:0]      o_icb_cmd_attri [SPLT_NUM-1:0];
    wire [SPLT_NUM-1:0] o_icb_rsp_valid;
    wire [SPLT_NUM-1:0] o_icb_rsp_ready;
    wire [SPLT_NUM-1:0] o_icb_rsp_err  ;
    wire [SPLT_NUM-1:0] o_icb_rsp_excl_ok  ;
    wire [DW-1:0] o_icb_rsp_rdata  [SPLT_NUM-1:0];
    wire [RSP_UW-1:0] o_icb_rsp_usr [SPLT_NUM-1:0];
    wire [SPLT_NUM-1:0] o_icb_cmd_ready_excpt_this [SPLT_NUM-1:0];
    wire sel_o_icb_cmd_ready;
    wire rspid_fifo_bypass;
    wire rspid_fifo_wen;
    wire rspid_fifo_ren;
    wire [SPLT_PTR_W-1:0] o_icb_rsp_port_id;
    wire rspid_fifo_i_valid;
    wire rspid_fifo_o_valid;
    wire rspid_fifo_o_valid_real;
    wire rspid_fifo_i_ready;
    wire rspid_fifo_i_ready_real;
    wire rspid_fifo_o_ready;
    wire [SPLT_FIFO_DW-1:0] rspid_fifo_rdat;
    wire [SPLT_FIFO_DW-1:0] rspid_fifo_rdat_real;
    wire [SPLT_FIFO_DW-1:0] rspid_fifo_wdat;
    wire rspid_fifo_full;
    reg [SPLT_PTR_W-1:0] i_splt_indic_id;
    wire i_icb_cmd_ready_pre;
    wire i_icb_cmd_valid_pre;
    wire i_icb_cmd_sel_pre;
    wire cmd_diff_branch_t[SPLT_NUM-1:0];
    wire i_icb_cmd_valid_pre2[SPLT_NUM-1:0];
    wire i_icb_cmd_sel_pre2[SPLT_NUM-1:0];
    wire i_icb_rsp_ready_pre;
    wire i_icb_rsp_valid_pre;
    for(i = 0; i < SPLT_NUM; i = i+1)
    begin:gen_icb_distract
      assign o_icb_cmd_ready[i]                             = o_bus_icb_cmd_ready[(i+1)*1     -1 : (i)*1     ];
      assign o_bus_icb_cmd_sel  [(i+1)*1     -1 : i*1     ] = o_icb_cmd_sel[i];
      assign o_bus_icb_cmd_valid[(i+1)*1     -1 : i*1     ] = o_icb_cmd_valid[i];
      assign o_bus_icb_cmd_read [(i+1)*1     -1 : i*1     ] = o_icb_cmd_read [i];
      assign o_bus_icb_cmd_addr [(i+1)*AW    -1 : i*AW    ] = o_icb_cmd_addr [i];
      assign o_bus_icb_cmd_wdata[(i+1)*DW    -1 : i*DW    ] = o_icb_cmd_wdata[i];
      assign o_bus_icb_cmd_wmask[(i+1)*DW/8    -1 : i*DW/8    ] = o_icb_cmd_wmask[i];
      assign o_bus_icb_cmd_beat [(i+1)*2     -1 : i*2     ] = o_icb_cmd_beat [i];
      assign o_bus_icb_cmd_lock [(i+1)*1     -1 : i*1     ] = o_icb_cmd_lock [i];
      assign o_bus_icb_cmd_excl [(i+1)*1     -1 : i*1     ] = o_icb_cmd_excl [i];
      assign o_bus_icb_cmd_size [(i+1)*3     -1 : i*3     ] = o_icb_cmd_size [i];
      assign o_bus_icb_cmd_usr  [(i+1)*CMD_UW -1 : i*CMD_UW ] = o_icb_cmd_usr  [i];
      assign o_bus_icb_cmd_xlen  [(i+1)*8 -1 : i*8 ] = o_icb_cmd_xlen  [i];
      assign o_bus_icb_cmd_xburst[(i+1)*2 -1 : i*2 ] = o_icb_cmd_xburst[i];
      assign o_bus_icb_cmd_modes [(i+1)*2 -1 : i*2 ] = o_icb_cmd_modes [i];
      assign o_bus_icb_cmd_dmode [(i+1)*1 -1 : i*1 ] = o_icb_cmd_dmode [i];
      assign o_bus_icb_cmd_attri [(i+1)*3 -1 : i*3 ] = o_icb_cmd_attri [i];
      assign o_bus_icb_rsp_ready[(i+1)*1-1 :i*1 ] = o_icb_rsp_ready[i];
      assign o_icb_rsp_valid[i]                   = o_bus_icb_rsp_valid[(i+1)*1-1 :i*1 ];
      assign o_icb_rsp_err  [i]                   = o_bus_icb_rsp_err  [(i+1)*1-1 :i*1 ];
      assign o_icb_rsp_excl_ok  [i]               = o_bus_icb_rsp_excl_ok  [(i+1)*1-1 :i*1 ];
      assign o_icb_rsp_rdata[i]                   = o_bus_icb_rsp_rdata[(i+1)*DW-1:i*DW];
      assign o_icb_rsp_usr       [i]              = o_bus_icb_rsp_usr  [(i+1)*RSP_UW-1:i*RSP_UW];
    end
    if(USE_ALL_READY == 1) begin:gen_all_ready
      assign sel_o_icb_cmd_ready = (&o_icb_cmd_ready);
    end
    else begin:gen_non_all_ready
      reg  sel_o_icb_cmd_ready_reg;
      always @ (*) begin : sel_o_icb_cmd_ready_PROC
        sel_o_icb_cmd_ready_reg = 1'b0;
          for(j = 0; j < SPLT_NUM; j = j+1) begin
            sel_o_icb_cmd_ready_reg = sel_o_icb_cmd_ready_reg | (i_icb_splt_indic_real[j] & o_icb_cmd_ready[j]);
          end
      end
      assign sel_o_icb_cmd_ready = sel_o_icb_cmd_ready_reg;
    end
    assign i_icb_cmd_ready_pre = sel_o_icb_cmd_ready;
    if(ALLOW_DIFF == 1) begin:gen_allow_diff
       assign i_icb_cmd_sel_pre       = i_icb_cmd_sel       & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre     = i_icb_cmd_valid     & (~rspid_fifo_full);
          for(i = 0; i < SPLT_NUM; i = i+1) begin:gen_allow_diff_splt_cmd
       assign cmd_diff_branch_t[i] = 1'b0;
       assign i_icb_cmd_sel_pre2  [i] = i_icb_cmd_sel       & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre2[i] = i_icb_cmd_valid     & (~rspid_fifo_full);
          end
       assign i_icb_cmd_ready     = i_icb_cmd_ready_pre & (~rspid_fifo_full);
    end
    else begin:gen_not_allow_diff
       wire cmd_diff_branch = (~rspid_fifo_empty) & (~(rspid_fifo_wdat[SPLT_PTR_W-1:0] == rspid_fifo_rdat_real[SPLT_PTR_W-1:0]));
       assign i_icb_cmd_sel_pre       = i_icb_cmd_sel       & (~cmd_diff_branch) & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre     = i_icb_cmd_valid     & (~cmd_diff_branch) & (~rspid_fifo_full);
        if(SPLT_PTR_1HOT == 1) begin:gen_pre2_ptr_1hot
          for(i = 0; i < SPLT_NUM; i = i+1) begin:gen_not_allow_diff_splt_cmd
       assign cmd_diff_branch_t[i] = (~rspid_fifo_empty) & (~(rspid_fifo_wdat[i] == rspid_fifo_rdat_real[i]));
       assign i_icb_cmd_sel_pre2   [i] = i_icb_cmd_sel       & (~cmd_diff_branch_t[i]) & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre2 [i] = i_icb_cmd_valid     & (~cmd_diff_branch_t[i]) & (~rspid_fifo_full);
          end
        end
        else begin: gen_pre2_ptr_not_1hot
          for(i = 0; i < SPLT_NUM; i = i+1) begin:gen_not_allow_diff_splt_cmd
       assign cmd_diff_branch_t[i] = 1'b0;
       assign i_icb_cmd_sel_pre2   [i] = i_icb_cmd_sel_pre;
       assign i_icb_cmd_valid_pre2 [i] = i_icb_cmd_valid_pre;
          end
        end
       assign i_icb_cmd_ready     = i_icb_cmd_ready_pre & (~cmd_diff_branch) & (~rspid_fifo_full);
    end
    if(SPLT_PTR_1HOT == 1) begin:gen_ptr_1hot
       always @ (*) begin : i_splt_indic_id_PROC
         i_splt_indic_id = i_icb_splt_indic_real;
       end
    end
    else begin:gen_ptr_not_1hot
       always @ (*) begin : i_splt_indic_id_PROC
         i_splt_indic_id = {SPLT_PTR_W{1'b0}};
         for(j = 0; j < SPLT_NUM; j = j+1) begin
// spyglass disable_block W216
// SMD: Inappropriate range select for int_part_sel variable
// SJ:  Here is not a real issue
           i_splt_indic_id = i_splt_indic_id | ({SPLT_PTR_W{i_icb_splt_indic_real[j]}} & (j[SPLT_PTR_W-1:0]));
// spyglass enable_block W216
         end
       end
    end
 if(ALLOW_DIFF == 1) begin:rspfifo_gen_allow_diff1
    assign rspid_fifo_wen = i_icb_cmd_valid & i_icb_cmd_ready;
    assign rspid_fifo_ren = i_icb_rsp_valid & i_icb_rsp_ready;
 end
 else begin: rspfifo_gen_allow_diff0
    assign rspid_fifo_wen = i_icb_cmd_valid & i_icb_cmd_ready 
                          ;
    assign rspid_fifo_ren = i_icb_rsp_valid & i_icb_rsp_ready 
                          ;
 end
    if(ALLOW_0CYCL_RSP == 1) begin: gen_allow_0rsp
        assign rspid_fifo_bypass = rspid_fifo_empty & rspid_fifo_wen & rspid_fifo_ren;
        assign o_icb_rsp_port_id = rspid_fifo_empty ? rspid_fifo_wdat[SPLT_PTR_W-1:0] : rspid_fifo_rdat_real[SPLT_PTR_W-1:0];
        assign i_icb_rsp_valid     = i_icb_rsp_valid_pre;
        assign i_icb_rsp_ready_pre = i_icb_rsp_ready;
    end
    else begin: gen_no_allow_0rsp
        assign rspid_fifo_bypass = 1'b0;
        assign o_icb_rsp_port_id = rspid_fifo_rdat_real[SPLT_PTR_W-1:0];
        assign i_icb_rsp_valid     = (~rspid_fifo_empty) & i_icb_rsp_valid_pre;
        assign i_icb_rsp_ready_pre = (~rspid_fifo_empty) & i_icb_rsp_ready;
    end
    assign rspid_fifo_i_valid = clk_en & rspid_fifo_wen & (~rspid_fifo_bypass);
    assign rspid_fifo_full    = (~rspid_fifo_i_ready_real);
    assign rspid_fifo_o_ready = clk_en & rspid_fifo_ren & (~rspid_fifo_bypass);
    assign rspid_fifo_empty   = (~rspid_fifo_o_valid_real);
      assign rspid_fifo_wdat   = i_splt_indic_id;
    assign rspid_fifo_o_valid_real = rspid_fifo_o_valid;
    assign rspid_fifo_i_ready_real = rspid_fifo_i_ready;
    assign rspid_fifo_rdat_real = rspid_fifo_rdat;
    if(FIFO_OUTS_NUM == 1) begin:gen_fifo_dp_1
      e603_subsys_gnrl_pipe_stage # (
        .CUT_READY (FIFO_CUT_READY),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (1),
        .DW  (SPLT_FIFO_DW)
      ) u_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else begin: gen_fifo_dp_gt_1
      e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT(FIFO_REG_OUT),
        .CUT_READY (FIFO_CUT_READY),
        .DP  (FIFO_OUTS_NUM),
        .DW  (SPLT_FIFO_DW)
      ) u_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    for(i = 0; i < SPLT_NUM; i = i+1)
    begin:gen_o_icb_cmd_valid
      for(ii = 0; ii < SPLT_NUM; ii = ii+1)
      begin:gen_o_cmd_ready_excpt_this
         if(i == ii) begin: gen_same_i
           assign o_icb_cmd_ready_excpt_this[i][ii] = 1'b1;
         end
         else begin: gen_no_same_i
           assign o_icb_cmd_ready_excpt_this[i][ii] = o_icb_cmd_ready[ii];
         end
      end
      if(USE_ALL_READY == 1) begin:gen_all_ready
         assign o_icb_cmd_valid[i] = i_icb_splt_indic_real[i] & i_icb_cmd_valid_pre2[i] & (&o_icb_cmd_ready_excpt_this[i]);
         assign o_icb_cmd_sel  [i] = i_icb_splt_indic_real[i] & i_icb_cmd_sel_pre2[i]   & (&o_icb_cmd_ready_excpt_this[i]);
      end
      else begin:gen_non_all_ready
         assign o_icb_cmd_valid[i] = i_icb_splt_indic_real[i] & i_icb_cmd_valid_pre2[i];
         assign o_icb_cmd_sel  [i] = i_icb_splt_indic_real[i] & i_icb_cmd_sel_pre2[i];
      end
      assign o_icb_cmd_lock[i] = i_icb_cmd_lock;
          assign o_icb_cmd_read [i] = i_icb_cmd_read ;
          assign o_icb_cmd_addr [i] = i_icb_cmd_addr ;
          assign o_icb_cmd_wdata[i] = i_icb_cmd_wdata;
          assign o_icb_cmd_wmask[i] = i_icb_cmd_wmask;
          assign o_icb_cmd_excl [i] = i_icb_cmd_excl ;
          assign o_icb_cmd_size [i] = i_icb_cmd_size ;
          assign o_icb_cmd_usr  [i] = i_icb_cmd_usr  ;
          assign o_icb_cmd_xburst[i] = i_icb_cmd_xburst;
          assign o_icb_cmd_modes [i] = i_icb_cmd_modes ;
          assign o_icb_cmd_dmode [i] = i_icb_cmd_dmode ;
          assign o_icb_cmd_attri [i] = i_icb_cmd_attri ;
          assign o_icb_cmd_xlen  [i] = i_icb_cmd_xlen  ;
          assign o_icb_cmd_beat [i] = i_icb_cmd_beat ;
    end
    if(SPLT_PTR_1HOT == 1) begin:gen_ptr_1hot_rsp
        for(i = 0; i < SPLT_NUM; i = i+1)
        begin:gen_o_icb_rsp_ready
          assign o_icb_rsp_ready[i] = (o_icb_rsp_port_id[i] & i_icb_rsp_ready_pre);
        end
        assign i_icb_rsp_valid_pre = |(o_icb_rsp_valid & o_icb_rsp_port_id);
        reg sel_i_icb_rsp_err;
        reg sel_i_icb_rsp_excl_ok;
        reg [DW-1:0] sel_i_icb_rsp_rdata;
        reg [RSP_UW-1:0] sel_i_icb_rsp_usr;
        always @ (*) begin : sel_icb_rsp_PROC
          sel_i_icb_rsp_err   = 1'b0;
          sel_i_icb_rsp_excl_ok   = 1'b0;
          sel_i_icb_rsp_rdata = {DW   {1'b0}};
          sel_i_icb_rsp_usr   = {RSP_UW{1'b0}};
          for(j = 0; j < SPLT_NUM; j = j+1) begin
            sel_i_icb_rsp_err     = sel_i_icb_rsp_err     | (       o_icb_rsp_port_id[j]   & o_icb_rsp_err[j]);
            sel_i_icb_rsp_excl_ok = sel_i_icb_rsp_excl_ok | (       o_icb_rsp_port_id[j]   & o_icb_rsp_excl_ok[j]);
            sel_i_icb_rsp_rdata   = sel_i_icb_rsp_rdata   | ({DW   {o_icb_rsp_port_id[j]}} & o_icb_rsp_rdata[j]);
            sel_i_icb_rsp_usr     = sel_i_icb_rsp_usr     | ({RSP_UW{o_icb_rsp_port_id[j]}} & o_icb_rsp_usr[j]);
          end
        end
        assign i_icb_rsp_err   = sel_i_icb_rsp_err  ;
        assign i_icb_rsp_excl_ok   = sel_i_icb_rsp_excl_ok  ;
        assign i_icb_rsp_rdata = sel_i_icb_rsp_rdata;
        assign i_icb_rsp_usr   = sel_i_icb_rsp_usr  ;
    end
    else begin:gen_ptr_not_1hot_rsp
        for(i = 0; i < SPLT_NUM; i = i+1)
        begin:gen_o_icb_rsp_ready
          assign o_icb_rsp_ready[i] = (o_icb_rsp_port_id == i[SPLT_PTR_W-1:0]) & i_icb_rsp_ready_pre;
        end
        assign i_icb_rsp_valid_pre = o_icb_rsp_valid[o_icb_rsp_port_id];
        assign i_icb_rsp_err     = o_icb_rsp_err    [o_icb_rsp_port_id];
        assign i_icb_rsp_excl_ok = o_icb_rsp_excl_ok[o_icb_rsp_port_id];
        assign i_icb_rsp_rdata   = o_icb_rsp_rdata  [o_icb_rsp_port_id];
        assign i_icb_rsp_usr     = o_icb_rsp_usr    [o_icb_rsp_port_id];
    end
  end
  endgenerate 
  assign splt_active = (i_icb_cmd_valid)
                     | (~rspid_fifo_empty)
                    ;
endmodule
module e603_subsys_gnrl_usr_ficb2ahbl
  #(
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter SUPPORT_LOCK = 0,
    parameter MON_DATA_WIDTH = 2,
    parameter AW = 32,
    parameter DW = 32
    )
  (
  input              icb_cmd_sel,
  input              icb_cmd_valid,
  output             icb_cmd_ready,
  input              icb_cmd_read,
  input  [AW-1:0]    icb_cmd_addr,
  input  [DW-1:0]    icb_cmd_wdata,
  input  [(DW/8-1):0]icb_cmd_wmask,
  input  [1:0]       icb_cmd_beat,
  input              icb_cmd_lock,
  input              icb_cmd_excl,
  input  [2:0]       icb_cmd_size,
  input  [7:0]       icb_cmd_xlen,
  input  [1:0]       icb_cmd_xburst,
  input  [1:0]       icb_cmd_modes,
  input              icb_cmd_dmode,
  input  [2:0]       icb_cmd_attri,
  input  [CMD_UW-1:0]    icb_cmd_usr,
  output [RSP_UW-1:0]    icb_rsp_usr,
  output [CMD_UW-1:0]    ahbl_huser,
  input  [RSP_UW-1:0]    ahbl_hruser,
  output             icb_rsp_valid,
  input              icb_rsp_ready,
  output             icb_rsp_err,
  output             icb_rsp_excl_ok,
  output [DW-1:0]    icb_rsp_rdata,
  output [1:0]       ahbl_htrans,
  output             ahbl_hwrite,
  output [AW    -1:0]ahbl_haddr,
  output [2:0]       ahbl_hsize,
  output             ahbl_hmastlock,
  output             ahbl_hexcl,
  output [2:0]       ahbl_hburst,
  output [DW    -1:0]ahbl_hwdata,
  output [3:0]       ahbl_hprot,
  output [1:0]       ahbl_hattri,
  output [1:0]       ahbl_master,
  input  [DW    -1:0]ahbl_hrdata,
  input  [1:0]       ahbl_hresp,
  input              ahbl_hresp_exok,
  input              ahbl_hready,
  input              bus_clk_en,
  output             icb2ahbl_pend_active,
  input              clk,
  input              rst_n
  );
  wire burst_flag_set;
  wire burst_flag_clr;
  wire burst_flag_r;
  wire             icb_cmd_read_r  ;
  wire [AW-1:0]    icb_cmd_addr_r  ;
  wire [DW-1:0]    icb_cmd_wdata_r ;
  wire [(DW/8-1):0]icb_cmd_wmask_r ;
  wire [2:0]       icb_cmd_size_r  ;
  wire [7:0]       icb_cmd_xlen_r  ;
  wire [1:0]       icb_cmd_xburst_r;
  wire [1:0]       icb_cmd_modes_r ;
  wire             icb_cmd_dmode_r ;
  wire [2:0]       icb_cmd_attri_r ;
  wire [CMD_UW-1:0]    icb_cmd_usr_r  ;
  wire            i_icb_rsp_valid;
  wire            i_icb_rsp_ready;
  wire            i_icb_rsp_err  ;
  wire            i_icb_rsp_excl_ok  ;
  wire [DW-1:0]   i_icb_rsp_rdata;
  wire [RSP_UW-1:0] i_icb_rsp_usr;
  localparam RSP_PACK_W = (2+DW
                           + RSP_UW
                     );
   e603_subsys_gnrl_dfflr #(1) icb_cmd_read_dfflr (burst_flag_set, icb_cmd_read, icb_cmd_read_r, clk, rst_n);// VPP_NO_REG_PARSE
   e603_subsys_gnrl_dfflr #(3) icb_cmd_size_dfflr (burst_flag_set, icb_cmd_size, icb_cmd_size_r, clk, rst_n);// VPP_NO_REG_PARSE
   e603_subsys_gnrl_dfflr #(8) icb_cmd_xlen_dfflr (burst_flag_set, icb_cmd_xlen, icb_cmd_xlen_r, clk, rst_n);// VPP_NO_REG_PARSE
   e603_subsys_gnrl_dfflr #(2) icb_cmd_xburst_dfflr (burst_flag_set, icb_cmd_xburst, icb_cmd_xburst_r, clk, rst_n);// VPP_NO_REG_PARSE
   e603_subsys_gnrl_dfflr #(2) icb_cmd_modes_dfflr (burst_flag_set, icb_cmd_modes, icb_cmd_modes_r, clk, rst_n);// VPP_NO_REG_PARSE
   e603_subsys_gnrl_dfflr #(1) icb_cmd_dmode_dfflr (burst_flag_set, icb_cmd_dmode, icb_cmd_dmode_r, clk, rst_n);// VPP_NO_REG_PARSE
   e603_subsys_gnrl_dfflr #(3) icb_cmd_attri_dfflr (burst_flag_set, icb_cmd_attri, icb_cmd_attri_r, clk, rst_n);// VPP_NO_REG_PARSE
   e603_subsys_gnrl_dfflr #(CMD_UW) icb_cmd_usr_dfflr (burst_flag_set, icb_cmd_usr, icb_cmd_usr_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire [1:0]        i_icb_cmd_xburst;
  wire [2:0]        i_icb_cmd_size;
  wire [7:0]        i_icb_cmd_xlen;
  wire i_icb_cmd_incr4 ;
  wire i_icb_cmd_incr8 ;
  wire i_icb_cmd_incr16;
  wire i_icb_cmd_incr4816;
  wire [AW-1:0] i_icb_cmd_addr_mask = ({AW{1'b1}} << i_icb_cmd_size);
  wire [AW-1:0] i_icb_cmd_addr_algned = (i_icb_cmd_addr_mask & ahbl_haddr);
  wire [10+1-1:0] i_icb_cmd_addr_incr =  (11'b1 << i_icb_cmd_size);
  wire [10+1 -1: 0] i_icb_cmd_addr_incr4816 = 
                     i_icb_cmd_incr4 ? (i_icb_cmd_addr_incr[10+1 -1: 0] << 2'd2) : 
                     i_icb_cmd_incr8 ? (i_icb_cmd_addr_incr[10+1 -1: 0] << 2'd3) : 
                                     (i_icb_cmd_addr_incr[10+1 -1: 0] << 3'd4) ;
// spyglass disable_block W484
// SMD: Possible loss of carry or borrow due to addition/subtraction
// SJ:  Here is not a real issue
  wire i_icb_cmd_addr_of;
  wire i_icb_cmd_addr_inc4816_of;
  wire [10-1:0] i_icb_cmd_addr_incr_size;
  wire [10-1:0] i_icb_cmd_addr_incr4816_size;
  assign {i_icb_cmd_addr_of, i_icb_cmd_addr_incr_size} = ({1'b0,i_icb_cmd_addr_algned[10-1:0]} + i_icb_cmd_addr_incr);
  assign {i_icb_cmd_addr_inc4816_of, i_icb_cmd_addr_incr4816_size} = ({1'b0,i_icb_cmd_addr_algned[10-1:0]} + i_icb_cmd_addr_incr4816
                                                                                                          - 1'd1);
  wire [10-1:0] i_icb_cmd_addr_wrap_mask = ((~{6'b0,i_icb_cmd_xlen[3:0]}) << i_icb_cmd_size);
  wire [10-1:0] i_icb_cmd_addr_incr_wrap = (i_icb_cmd_addr_incr_size & (~i_icb_cmd_addr_wrap_mask)) 
                                       | (ahbl_haddr[10-1:0] & i_icb_cmd_addr_wrap_mask);
// spyglass enable_block W484
  wire i_icb_cmd_fxed = (i_icb_cmd_xburst == 2'b00);
  wire i_icb_cmd_wrap = (i_icb_cmd_xburst == 2'b10);
  wire [AW-1:0] i_icb_cmd_addr_nxt = i_icb_cmd_fxed ? ahbl_haddr : 
                                 i_icb_cmd_wrap ? {ahbl_haddr[AW-1:10],i_icb_cmd_addr_incr_wrap} :
                                                 {ahbl_haddr[AW-1:10],i_icb_cmd_addr_incr_size};
  wire burst_valid_r;
  wire burst_valid_real;
  wire ahbl_eff_trans;
 wire [AW-1:0] icb_cmd_addr_ofst;
 wire icb_cmd_addr_ena = (burst_flag_set | ((~burst_flag_clr) & burst_flag_r & icb_cmd_valid & icb_cmd_ready)) & bus_clk_en;
e603_subsys_gnrl_dfflr #(AW) icb_cmd_addr_dfflr (icb_cmd_addr_ena, i_icb_cmd_addr_nxt, icb_cmd_addr_r, clk, rst_n);// VPP_NO_REG_PARSE
 wire icb_cmd_valid_msked;
 wire i_icb_cmd_incr_no4816;
 wire icb_cmd_incr_no4816_1stovf = i_icb_cmd_incr_no4816 & icb_cmd_valid_msked & icb_cmd_beat[0] & i_icb_cmd_addr_of;
  wire cmd_sel_r = ((~icb_cmd_valid) & burst_flag_r);
  wire              i_icb_cmd_read   = cmd_sel_r ? icb_cmd_read_r   : icb_cmd_read  ;
  wire [AW-1:0]     i_icb_cmd_addr   = cmd_sel_r ? icb_cmd_addr_r   : icb_cmd_addr  ;
  wire [CMD_UW-1:0] i_icb_cmd_usr   = cmd_sel_r ? icb_cmd_usr_r   : icb_cmd_usr  ;
  assign            i_icb_cmd_size   = cmd_sel_r ? icb_cmd_size_r   : icb_cmd_size  ;
  assign            i_icb_cmd_xlen   = cmd_sel_r ? icb_cmd_xlen_r   : icb_cmd_xlen  ;
  assign            i_icb_cmd_xburst = cmd_sel_r ? icb_cmd_xburst_r : icb_cmd_xburst;
  wire [1:0]        i_icb_cmd_modes  = cmd_sel_r ? icb_cmd_modes_r  : icb_cmd_modes ;
  wire              i_icb_cmd_dmode  = cmd_sel_r ? icb_cmd_dmode_r  : icb_cmd_dmode ;
  wire [2:0]        i_icb_cmd_attri  = cmd_sel_r ? icb_cmd_attri_r  : icb_cmd_attri ;
 wire icb_cmd_hsked;
 wire i_icb_cmd_hsked;
 assign i_icb_cmd_hsked = icb_cmd_hsked;
 wire i_icb_cmd_beat_end = icb_cmd_beat[1];
 wire icb_cmd_1kend_r;
 wire icb_cmd_1kend_set = (
                            i_icb_cmd_hsked
                            ) & (
                             icb_cmd_incr_no4816_1stovf |
                             (burst_flag_r 
                                     & (~i_icb_cmd_beat_end)
                                     & i_icb_cmd_incr_no4816 & i_icb_cmd_addr_of)
                             );
 wire icb_cmd_1kend_clr = i_icb_cmd_hsked & icb_cmd_1kend_r;
 wire icb_cmd_1kend_ena = (icb_cmd_1kend_set | icb_cmd_1kend_clr) & bus_clk_en;
 wire icb_cmd_1kend_nxt = ~icb_cmd_1kend_clr;
e603_subsys_gnrl_dfflr #(1) icb_cmd_1kend_dfflr (icb_cmd_1kend_ena, icb_cmd_1kend_nxt, icb_cmd_1kend_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_cmd_incr4816_of = (icb_cmd_valid_msked & icb_cmd_beat[0] & i_icb_cmd_incr4816 & i_icb_cmd_addr_inc4816_of);
  wire ahbl_hready_en = ahbl_hready & bus_clk_en;
  wire lock2idle_r;
  wire lock_flag_r;
  assign ahbl_eff_trans = ahbl_hready_en & ahbl_htrans[1];
  assign icb_cmd_hsked = icb_cmd_valid & icb_cmd_ready;
 assign burst_flag_set = ((icb_cmd_beat[0] & icb_cmd_hsked 
                                    & (~icb_cmd_incr_no4816_1stovf)
                                    & (~icb_cmd_incr4816_of)
                                    ) 
                                    | (icb_cmd_1kend_clr & (~i_icb_cmd_beat_end))
                                    ) 
                      & (ahbl_hburst != 3'b000);
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 i_icb_rsp_err,
                                 i_icb_rsp_excl_ok,
                                 i_icb_rsp_rdata 
                                ,i_icb_rsp_usr
                                 };
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 icb_rsp_err,
                                 icb_rsp_excl_ok,
                                 icb_rsp_rdata 
                                ,icb_rsp_usr
                                 } = rsp_fifo_o_dat;
    assign icb_rsp_valid   = i_icb_rsp_valid; 
    assign i_icb_rsp_ready = icb_rsp_ready; 
    assign rsp_fifo_o_dat = rsp_fifo_i_dat;
    wire i_icb_rsp_fifo_avail = 1'b1;
 assign burst_flag_clr = ((icb_cmd_beat[1] & icb_cmd_hsked) | icb_cmd_1kend_set) & burst_flag_r;
 assign burst_valid_r = 1'b0;
 assign burst_valid_real = 1'b0;
 wire burst_flag_ena = (burst_flag_set |   burst_flag_clr) & bus_clk_en;
 wire burst_flag_nxt = (~burst_flag_clr);
e603_subsys_gnrl_dfflr #(1) burst_flag_dfflr (burst_flag_ena, burst_flag_nxt, burst_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_cmd_ready  = ahbl_hready_en   & (~lock2idle_r) & i_icb_rsp_fifo_avail & (~burst_valid_r);
  assign ahbl_htrans[1] = (icb_cmd_valid_msked | burst_valid_real) & (~lock2idle_r);
  assign ahbl_htrans[0] = burst_flag_r;
  assign icb_cmd_valid_msked = (icb_cmd_valid & i_icb_rsp_fifo_avail & (~burst_valid_r));
  localparam FSM_W  = 2;
  localparam STA_AR = 2'b00;
  localparam STA_WD = 2'b01;
  localparam STA_RD = 2'b10;
  wire[FSM_W-1:0] ahbl_sta_r;
  wire[FSM_W-1:0] ahbl_sta_nxt;
  wire to_wd_sta = ahbl_eff_trans & ahbl_hwrite;
  wire to_rd_sta = ahbl_eff_trans & (~ahbl_hwrite);
  wire to_ar_sta = ahbl_hready_en & (~ahbl_htrans[1]);
  wire  ahbl_sta_is_ar = (ahbl_sta_r == STA_AR);
  assign ahbl_sta_nxt = ahbl_hready_en ?  (
                               {FSM_W{to_ar_sta}} & (STA_AR)
                             | {FSM_W{to_wd_sta}} & (STA_WD)
                             | {FSM_W{to_rd_sta}} & (STA_RD)
                         ) : ahbl_sta_r;
e603_subsys_gnrl_dffr #(FSM_W) ahbl_sta_dffr (ahbl_sta_nxt, ahbl_sta_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire [DW-1:0]ahbl_hwdata_r;
  wire ahbl_hwdata_ena = to_wd_sta;
e603_subsys_gnrl_dfflr #(DW) ahbl_hwdata_dfflr (ahbl_hwdata_ena, icb_cmd_wdata, ahbl_hwdata_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign ahbl_hwrite = ~i_icb_cmd_read;
  assign ahbl_haddr  = i_icb_cmd_addr;
  assign ahbl_huser  = i_icb_cmd_usr;
  assign ahbl_hsize  = i_icb_cmd_size;
  assign ahbl_hexcl  = 1'b0;
  wire icb_cmd_burst_fixd = (i_icb_cmd_xburst == 2'b00);
  wire i_icb_cmd_burst_incr = (i_icb_cmd_xburst == 2'b01);
  wire icb_cmd_burst_wrap = (i_icb_cmd_xburst == 2'b10);
  wire icb_cmd_xlen_0  = (i_icb_cmd_xlen == 8'd0);
  wire icb_cmd_xlen_4  = (i_icb_cmd_xlen == 8'd3);
  wire icb_cmd_xlen_8  = (i_icb_cmd_xlen == 8'd7);
  wire icb_cmd_xlen_16 = (i_icb_cmd_xlen == 8'd15);
  wire icb_cmd_wrap4 = icb_cmd_burst_wrap & icb_cmd_xlen_4;
  wire icb_cmd_wrap8 = icb_cmd_burst_wrap & icb_cmd_xlen_8;
  wire icb_cmd_wrap16 = icb_cmd_burst_wrap & icb_cmd_xlen_16;
  assign i_icb_cmd_incr4 = i_icb_cmd_burst_incr & icb_cmd_xlen_4;
  assign i_icb_cmd_incr8 = i_icb_cmd_burst_incr & icb_cmd_xlen_8;
  assign i_icb_cmd_incr16 = i_icb_cmd_burst_incr & icb_cmd_xlen_16;
  assign i_icb_cmd_incr4816 = i_icb_cmd_incr4 | i_icb_cmd_incr8 | i_icb_cmd_incr16;
  assign i_icb_cmd_incr_no4816 = i_icb_cmd_burst_incr & (~i_icb_cmd_incr4816);
  wire ahbl_is_burst = (icb_cmd_valid_msked & icb_cmd_beat[0]) | burst_flag_r;
  assign ahbl_hburst = (icb_cmd_incr4816_of | icb_cmd_incr_no4816_1stovf) ? 3'b000 : 
                       (ahbl_is_burst & icb_cmd_wrap4) ? 3'b010 :
                       (ahbl_is_burst & i_icb_cmd_incr4) ? 3'b011 :
                       (ahbl_is_burst & icb_cmd_wrap8) ? 3'b100 :
                       (ahbl_is_burst & i_icb_cmd_incr8) ? 3'b101 :
                       (ahbl_is_burst & icb_cmd_wrap16) ? 3'b110 :
                       (ahbl_is_burst & i_icb_cmd_incr16) ? 3'b111 :
                       (ahbl_is_burst & (i_icb_cmd_burst_incr & (~icb_cmd_xlen_0))) ? 3'b001 : 3'b000;
  assign ahbl_hwdata = ahbl_hwdata_r;
  wire icb_cmd_mmode  = (i_icb_cmd_modes == 2'd0);
  wire icb_cmd_hmode  = (i_icb_cmd_modes == 2'd1);
  wire icb_cmd_smode  = (i_icb_cmd_modes == 2'd2);
  wire icb_cmd_umode  = (i_icb_cmd_modes == 2'd3);
  wire icb_cmd_ifu    = i_icb_cmd_attri[0];
  wire icb_cmd_device = (~(i_icb_cmd_attri[2] & i_icb_cmd_attri[1])) & i_icb_cmd_attri[1];
  wire icb_cmd_nc     = (~(i_icb_cmd_attri[2] & i_icb_cmd_attri[1])) & i_icb_cmd_attri[2];
  assign ahbl_hprot[0] = (~icb_cmd_ifu);
  assign ahbl_hprot[1] = icb_cmd_mmode;
  assign ahbl_hprot[2] = (~icb_cmd_device); 
  assign ahbl_hprot[3] = (~icb_cmd_device) & (~icb_cmd_nc);
  assign ahbl_hattri = (icb_cmd_nc | icb_cmd_device) ? 2'b00 : 2'b11;
  wire icb_cmd_from_ifu  = (~i_icb_cmd_dmode) & (~ahbl_hprot[0]);
  wire icb_cmd_from_data = (~i_icb_cmd_dmode) & ahbl_hprot[0];
  wire icb_cmd_from_dbg  = i_icb_cmd_dmode;
  wire [1:0] icb_cmd_master =
                        icb_cmd_from_data ? 2'b00 :
                        icb_cmd_from_dbg ? 2'b01 :
                        icb_cmd_from_ifu ? 2'b10 :
                                      2'b11;
  assign ahbl_master = icb_cmd_master;
  assign i_icb_rsp_valid = ahbl_hready & (~ahbl_sta_is_ar);
  assign i_icb_rsp_rdata = ahbl_hrdata;
  assign i_icb_rsp_usr = ahbl_hruser;
  assign i_icb_rsp_err   = ahbl_hresp[0];
  assign i_icb_rsp_excl_ok   = ahbl_hresp_exok;
  wire lock2idle_set;
  wire lock2idle_clr;
  wire lock2idle_ena;
  wire lock2idle_nxt;
  wire lock_flag_set;
  wire lock_flag_clr;
  wire lock_flag_ena;
  wire lock_flag_nxt;
  generate
    if(SUPPORT_LOCK == 1) begin:gen_lock_1
      assign ahbl_hmastlock    = ((icb_cmd_lock & icb_cmd_valid) | lock_flag_r)
                           & (~lock2idle_r)  
                           & (~(
                                  ((~icb_cmd_lock) & icb_cmd_valid)
                               )
                             );
      assign lock2idle_set = lock_flag_clr;
      assign lock2idle_clr = lock2idle_r & to_ar_sta;
      assign lock2idle_ena = (lock2idle_set | lock2idle_clr) & bus_clk_en;
      assign lock2idle_nxt = lock2idle_set & (~lock2idle_clr);
e603_subsys_gnrl_dfflr #(1) lock2idle_dfflr (lock2idle_ena, lock2idle_nxt, lock2idle_r, clk, rst_n);// VPP_NO_REG_PARSE
      assign lock_flag_set = (ahbl_eff_trans & icb_cmd_lock);
      assign lock_flag_clr = lock_flag_r & (
                             (ahbl_eff_trans & (~icb_cmd_lock))
                           )
                           ;
      assign lock_flag_ena = (lock_flag_set | lock_flag_clr) & bus_clk_en;
      assign lock_flag_nxt = lock_flag_set & (~lock_flag_clr);
e603_subsys_gnrl_dfflr #(1) lock_flag_dfflr (lock_flag_ena, lock_flag_nxt, lock_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
    end
    else begin: gen_lock_0
      assign lock2idle_set = 1'b0;
      assign lock2idle_clr = 1'b0;
      assign lock2idle_ena = 1'b0;
      assign lock2idle_nxt = 1'b0;
      assign lock_flag_set = 1'b0;
      assign lock_flag_clr = 1'b0;
      assign lock_flag_ena = 1'b0;
      assign lock_flag_nxt = 1'b0;
      assign ahbl_hmastlock= 1'b0;
      assign lock2idle_r   = 1'b0;
      assign lock_flag_r   = 1'b0;
    end
  endgenerate
  assign icb2ahbl_pend_active = lock2idle_r;
endmodule
module e603_subsys_gnrl_usr_ahbl2ficb
  #(
    parameter OUTS_CNT_W = 2,
    parameter SUPPORT_ICB_BURST = 0,
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter WR_EARLY_RETURN = 1,
    parameter AW = 32,
    parameter DW = 32  
    )
  (
  input              bus_clk_en,
  output             ahbl2icb_active,
  output  [RSP_UW-1:0] ahbl_hruser,
  input  [RSP_UW-1:0]  icb_rsp_usr,
  input              ahbl_hsel,
  input              ahbl_hexcl,
  input  [1:0]       ahbl_htrans,
  input              ahbl_hwrite,
  input  [AW    -1:0]ahbl_haddr,
  input  [2:0]       ahbl_hsize,
  input  [3:0]       ahbl_hprot,
  input  [DW    -1:0]ahbl_hwdata,
  input  [CMD_UW-1:0]    ahbl_huser,
  input              ahbl_hmastlock,
  input  [2:0]       ahbl_hburst,
  output  [DW   -1:0]ahbl_hrdata,
  output  [1:0]      ahbl_hresp,
  output             ahbl_hresp_exok,
  input              ahbl_hready_in,
  output             ahbl_hready_out,
  output             icb_cmd_sel,
  output             icb_cmd_valid,
  input              icb_cmd_ready,
  output             icb_cmd_read,
  output  [AW-1:0]   icb_cmd_addr,
  output  [CMD_UW-1:0]   icb_cmd_usr,
  output  [DW-1:0]   icb_cmd_wdata,
  output  [(DW/8-1):0] icb_cmd_wmask,
  output  [2:0]      icb_cmd_size,
  output             icb_cmd_excl,
  output             icb_cmd_lock,
  output [7:0]       icb_cmd_xlen,
  output [1:0]       icb_cmd_beat,
  output [1:0]       icb_cmd_xburst,
  output [1:0]       icb_cmd_modes,
  output             icb_cmd_dmode,
  output [2:0]       icb_cmd_attri,
  input              icb_rsp_valid, 
  output             icb_rsp_ready,
  input              icb_rsp_err,
  input              icb_rsp_excl_ok,
  input  [DW-1:0]    icb_rsp_rdata,
  input              clk,
  input              rst_n
  );
  wire ahbl_hmastlock_r;
  wire  i_icb_cmd_valid;
  wire  i_icb_cmd_ready;
  wire  i_icb_cmd_read;
  wire  i_icb_cmd_excl;
  wire  [AW-1:0] i_icb_cmd_addr;
  wire  [CMD_UW-1:0] i_icb_cmd_usr;
  wire  [DW-1:0] i_icb_cmd_wdata;
  wire  [(DW/8-1):0] i_icb_cmd_wmask;
  wire  [3-1:0] i_icb_cmd_size;
  wire        i_icb_cmd_lock;
  wire [7:0] i_icb_cmd_xlen;
  wire [1:0] i_icb_cmd_xburst;
  wire [1:0] i_icb_cmd_beat;
  wire [1:0] i_icb_cmd_modes;
  wire       i_icb_cmd_dmode;
  wire [2:0] i_icb_cmd_attri;
  localparam BUF_CMD_PACK_W = (AW+DW+(DW/8)+5+1+1+8+2+2+CMD_UW+3+2) 
        ;
  wire [BUF_CMD_PACK_W-1:0] icb_cmd_pack;
  wire [BUF_CMD_PACK_W-1:0] i_icb_cmd_pack =  {
                      i_icb_cmd_read,
                      i_icb_cmd_excl,
                      i_icb_cmd_addr,
                      i_icb_cmd_usr,
                      i_icb_cmd_wdata,
                      i_icb_cmd_wmask,
                      i_icb_cmd_size,
                      i_icb_cmd_lock,
                     i_icb_cmd_xlen,
                     i_icb_cmd_xburst,
                     i_icb_cmd_beat,
                     i_icb_cmd_modes,
                     i_icb_cmd_dmode,
                     i_icb_cmd_attri 
                    };
  assign {
                      icb_cmd_read,
                      icb_cmd_excl,
                      icb_cmd_addr,
                                          icb_cmd_usr,
                      icb_cmd_wdata,
                      icb_cmd_wmask,
                      icb_cmd_size,
                      icb_cmd_lock,
                     icb_cmd_xlen,
                     icb_cmd_xburst,
                     icb_cmd_beat,
                     icb_cmd_modes,
                     icb_cmd_dmode,
                     icb_cmd_attri 
                    } = icb_cmd_pack;
  wire cmd_bypbuf_fifo_o_vld;
  wire outs_cnt_max;
  wire i_icb_cmd_valid_raw;
  wire i_icb_cmd_ready_raw;
  assign i_icb_cmd_valid_raw = i_icb_cmd_valid     & (~outs_cnt_max);
  assign i_icb_cmd_ready     = i_icb_cmd_ready_raw & (~outs_cnt_max);
  e603_subsys_gnrl_bypbuf # (
   .DP(1),
   .DW(BUF_CMD_PACK_W)
  ) u_byp_icb_cmd_buf(
    .i_vld(i_icb_cmd_valid_raw & bus_clk_en),
    .i_rdy(i_icb_cmd_ready_raw),
    .i_dat(i_icb_cmd_pack),
    .o_vld(icb_cmd_valid),
    .o_rdy(icb_cmd_ready & bus_clk_en),
    .o_dat(icb_cmd_pack),
    .fifo_o_vld(cmd_bypbuf_fifo_o_vld),
    .clk  (clk  ),
    .rst_n(rst_n)
   );
  wire i_icb_rsp_valid_raw;
  wire i_icb_rsp_ready_raw;
  wire i_icb_rsp_valid;
  wire i_icb_rsp_ready;
  wire i_icb_rsp_err;
  wire i_icb_rsp_excl_ok;
  wire [DW-1:0] i_icb_rsp_rdata;
  wire [RSP_UW-1:0] i_icb_rsp_usr;
  localparam BUF_RSP_PACK_W = (DW+2) 
            + RSP_UW
        ;
  wire [BUF_RSP_PACK_W-1:0]i_icb_rsp_pack;
  wire [BUF_RSP_PACK_W-1:0]icb_rsp_pack;
  assign icb_rsp_pack = {
                          icb_rsp_excl_ok,
                          icb_rsp_err,
                          icb_rsp_usr,
                          icb_rsp_rdata
                          };
  assign {
                          i_icb_rsp_excl_ok,
                          i_icb_rsp_err,
                          i_icb_rsp_usr,
                          i_icb_rsp_rdata
                          } = i_icb_rsp_pack;
  e603_subsys_gnrl_bypbuf # (
    .DP(1),
    .DW(BUF_RSP_PACK_W)
  ) u_rsp_bypbuf(
      .i_vld   (icb_rsp_valid & bus_clk_en),
      .i_rdy   (icb_rsp_ready),
      .o_vld   (i_icb_rsp_valid_raw),
      .o_rdy   (i_icb_rsp_ready_raw & bus_clk_en),
      .i_dat   (icb_rsp_pack),
      .o_dat   (i_icb_rsp_pack),
      .fifo_o_vld(),
      .clk     (clk  ),
      .rst_n   (rst_n)
  );
  wire ahbl_hready_real = ahbl_hready_out & ahbl_hready_in & bus_clk_en;
  wire ahbl_hsel_trans_busy  =
        ahbl_hsel
      & ahbl_htrans[0]
      ;
  wire ahbl_hsel_trans  =
        ahbl_hsel
      & ahbl_htrans[1]
      ;
  wire ahbl_addr_en  = ahbl_hsel_trans
      & ahbl_hready_real;
  wire [1:0] ahbl_htrans_r;
  wire ahbl_data_en  =
        ahbl_htrans_r[1]
      & ahbl_hready_real;
  wire ahbl_hvalid_r;
  wire ahbl_hvalid_ena = ahbl_hready_real;
  wire ahbl_hvalid_nxt = ahbl_addr_en;
e603_subsys_gnrl_dfflr #(1) ahbl_hvalid_dfflr (ahbl_hvalid_ena, ahbl_hvalid_nxt, ahbl_hvalid_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_htrans_ena = ahbl_hready_real;
  wire [1:0] ahbl_htrans_nxt = ahbl_htrans;
e603_subsys_gnrl_dfflr #(2) ahbl_htrans_dfflr (ahbl_htrans_ena, ahbl_htrans_nxt, ahbl_htrans_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_hexcl_tie = 1'b0;
  wire ahbl_hexcl_r;
  wire ahbl_hexcl_ena = ahbl_hready_real;
  wire ahbl_hexcl_nxt = ahbl_hexcl_tie;
e603_subsys_gnrl_dfflr #(1) ahbl_hexcl_dfflr (ahbl_hexcl_ena, ahbl_hexcl_nxt, ahbl_hexcl_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_hwrite_r;
  wire ahbl_hwrite_ena = ahbl_hready_real;
  wire ahbl_hwrite_nxt = ahbl_hwrite;
e603_subsys_gnrl_dfflr #(1) ahbl_hwrite_dfflr (ahbl_hwrite_ena, ahbl_hwrite_nxt, ahbl_hwrite_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_hmastlock_ena = ahbl_hready_real;
  wire ahbl_hmastlock_nxt = 
                         ahbl_hmastlock;
e603_subsys_gnrl_dfflr #(1) ahbl_hmastlock_dfflr (ahbl_hmastlock_ena, ahbl_hmastlock_nxt, ahbl_hmastlock_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire [2:0] ahbl_hburst_r;
  wire ahbl_hburst_ena = ahbl_hready_real;
  wire [2:0] ahbl_hburst_nxt = ahbl_hburst[2:0];
e603_subsys_gnrl_dfflr #(3) ahbl_hburst_dfflr (ahbl_hburst_ena, ahbl_hburst_nxt, ahbl_hburst_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire [2:0] ahbl_hsize_r;
  wire ahbl_hsize_ena = ahbl_hready_real;
  wire [2:0] ahbl_hsize_nxt = ahbl_hsize[2:0];
e603_subsys_gnrl_dfflr #(3) ahbl_hsize_dfflr (ahbl_hsize_ena, ahbl_hsize_nxt, ahbl_hsize_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_haddr_ena = ahbl_hready_real;
  wire [AW-1:0] ahbl_haddr_r;
  wire [AW-1:0] ahbl_haddr_nxt = ahbl_haddr;
e603_subsys_gnrl_dfflr #(AW) ahbl_haddr_dfflr (ahbl_haddr_ena, ahbl_haddr_nxt, ahbl_haddr_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_huser_ena = ahbl_hready_real;
  wire [CMD_UW-1:0] ahbl_huser_r;
  wire [CMD_UW-1:0] ahbl_huser_nxt = ahbl_huser;
e603_subsys_gnrl_dfflr #(CMD_UW) ahbl_huser_dfflr (ahbl_huser_ena, ahbl_huser_nxt, ahbl_huser_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_hprot_ena = ahbl_hready_real;
  wire [3:0] ahbl_hprot_r;
  wire [3:0] ahbl_hprot_nxt = ahbl_hprot;
e603_subsys_gnrl_dfflr #(4) ahbl_hprot_dfflr (ahbl_hprot_ena, ahbl_hprot_nxt, ahbl_hprot_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_wr_vld_r;
  wire[3-1:0] i_icb_cmd_burst = icb_wr_vld_r ? ahbl_hburst_r[2:0] : ahbl_hburst[2:0];
  assign i_icb_cmd_read = icb_wr_vld_r ? (~ahbl_hwrite_r) : (~ahbl_hwrite);
  assign i_icb_cmd_addr = icb_wr_vld_r ? ahbl_haddr_r : ahbl_haddr;
  assign i_icb_cmd_usr  = icb_wr_vld_r ? ahbl_huser_r : ahbl_huser;
  assign i_icb_cmd_size = icb_wr_vld_r ? ahbl_hsize_r : ahbl_hsize;
  assign i_icb_cmd_lock = 1'b0;
  assign i_icb_cmd_excl = 1'b0;
  assign i_icb_cmd_wdata = ahbl_hwdata;
  generate
  if(SUPPORT_ICB_BURST == 1) begin: icb_burst_gen
      assign i_icb_cmd_xlen   =
                      ((i_icb_cmd_burst == 3'b010) | (i_icb_cmd_burst == 3'b011)) ? 8'd3 :
                      ((i_icb_cmd_burst == 3'b100) | (i_icb_cmd_burst == 3'b101)) ? 8'd7 :
                      ((i_icb_cmd_burst == 3'b110) | (i_icb_cmd_burst == 3'b111)) ? 8'd15 : 8'd0;
      assign i_icb_cmd_xburst =
                           ((i_icb_cmd_burst == 3'b010) | (i_icb_cmd_burst == 3'b100) | (i_icb_cmd_burst == 3'b110)) ? 2'b10 : 
                           ((i_icb_cmd_burst == 3'b011) | (i_icb_cmd_burst == 3'b101) | (i_icb_cmd_burst == 3'b111)) ? 2'b01 : 
                           2'b0;
      wire       burst_last;
      wire [3:0] burst_cnt_r;
      wire [3:0] burst_cnt_nxt;
      wire       burst_cnt_ena;
      wire burst_trans = (i_icb_cmd_xburst != 2'b0);
      wire burst_first = (burst_cnt_r == 4'd0);
      assign burst_cnt_nxt = burst_last ? 4'b0 : (burst_cnt_r + 4'b1);
      assign burst_last = (burst_cnt_r == i_icb_cmd_xlen[3:0]) & (~burst_first);
      assign burst_cnt_ena = (i_icb_cmd_xburst !=2'b0) & i_icb_cmd_valid && i_icb_cmd_ready & bus_clk_en;
e603_subsys_gnrl_dfflr #(4) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
      assign i_icb_cmd_beat[0] = burst_first & burst_trans;
      assign i_icb_cmd_beat[1] = burst_last  & burst_trans;
  end
  else begin: no_icb_burst_gen
      assign i_icb_cmd_xlen   = 8'd0;
      assign i_icb_cmd_xburst = 2'b0;
      assign i_icb_cmd_beat[0] = 1'b0;
      assign i_icb_cmd_beat[1] = 1'b0;
  end
  endgenerate
  wire i_icb_cmd_mmode = icb_wr_vld_r ? (ahbl_hprot_r[1]) : (ahbl_hprot[1]);
  assign i_icb_cmd_modes = i_icb_cmd_mmode ? 2'd0 : 2'd3; 
  assign i_icb_cmd_dmode = 1'b0;
  assign i_icb_cmd_attri[0] = icb_wr_vld_r ? (~ahbl_hprot_r[0]) : (~ahbl_hprot[0]);
  assign i_icb_cmd_attri[1] = icb_wr_vld_r ? (~ahbl_hprot_r[2]) : (~ahbl_hprot[2]);
  assign i_icb_cmd_attri[2] = icb_wr_vld_r ? (~ahbl_hprot_r[3] & ahbl_hprot_r[2]) : (~ahbl_hprot[3] & ahbl_hprot[2]);
  wire ahbl_hwrite_device = (~ahbl_hprot[2]);
  wire [(DW/8-1):0] ahbl2icb_wmask;
  wire [(DW/8-1):0] ahbl2icb_wmask_r;
  wire ahbl2icb_wmask_ena = ahbl_hready_real;
  wire [(DW/8-1):0] ahbl2icb_wmask_nxt = ahbl2icb_wmask;
e603_subsys_gnrl_dfflr #(DW/8) ahbl2icb_wmask_dfflr (ahbl2icb_wmask_ena, ahbl2icb_wmask_nxt, ahbl2icb_wmask_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign i_icb_cmd_wmask = ahbl2icb_wmask_r;
  generate
  if(DW == 64) begin:gen_dw_64
     assign ahbl2icb_wmask =
         (ahbl_hsize == 3'b00) ? (1'b1 << ahbl_haddr[2:0])
       : (ahbl_hsize == 3'b01) ? (2'b11 << {ahbl_haddr[2:1],1'b0})
       : (ahbl_hsize == 3'b10) ? (4'b1111 << {ahbl_haddr[2],2'b0})
       : (8'b1111_1111)
       ;
  end
  if(DW == 32) begin:gen_dw_32
     assign ahbl2icb_wmask =
         (ahbl_hsize == 3'b00) ? (1'b1 << ahbl_haddr[1:0])
       : (ahbl_hsize == 3'b01) ? (2'b11 << {ahbl_haddr[1:1],1'b0})
       : (ahbl_hsize == 3'b10) ? (4'b1111)
       : (4'b1111)
       ;
  end
  endgenerate
  wire rd_hresp_1st_err_r;
  wire rd_hresp_1st_err;
  wire rd_hresp_1st_err_set = i_icb_rsp_valid & rd_hresp_1st_err  & bus_clk_en;
  wire rd_hresp_1st_err_clr = rd_hresp_1st_err_r & ahbl_hready_real;
  wire rd_hresp_1st_err_ena = rd_hresp_1st_err_set | rd_hresp_1st_err_clr;
  wire rd_hresp_1st_err_nxt = rd_hresp_1st_err_set | (~rd_hresp_1st_err_clr);
e603_subsys_gnrl_dfflr #(1) rd_hresp_1st_err_dfflr (rd_hresp_1st_err_ena, rd_hresp_1st_err_nxt, rd_hresp_1st_err_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_hsel_trans_wr = (ahbl_hsel_trans & ahbl_hwrite);
  wire icb_wr_vld_set = ahbl_hvalid_ena & ahbl_hsel_trans_wr & bus_clk_en;
  wire icb_wr_vld_clr = i_icb_cmd_valid & i_icb_cmd_ready & (~i_icb_cmd_read) & bus_clk_en;
  wire icb_wr_vld_ena = icb_wr_vld_set | icb_wr_vld_clr;
  wire icb_wr_vld_nxt = icb_wr_vld_set | (~icb_wr_vld_clr);
e603_subsys_gnrl_dfflr #(1) icb_wr_vld_dfflr (icb_wr_vld_ena, icb_wr_vld_nxt, icb_wr_vld_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_hwrite_device_r;
  wire ahbl_hwrite_device_set = icb_wr_vld_set;
  wire ahbl_hwrite_device_clr = icb_wr_vld_clr;
  wire ahbl_hwrite_device_ena = ahbl_hwrite_device_set | ahbl_hwrite_device_clr;
  wire ahbl_hwrite_device_nxt = ahbl_hwrite_device_set ? ahbl_hwrite_device : 1'b0;
e603_subsys_gnrl_dfflr #(1) ahbl_hwrite_device_dfflr                (ahbl_hwrite_device_ena, ahbl_hwrite_device_nxt, ahbl_hwrite_device_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_noearly_vld_r;
  wire icb_noearly_vld_set;
  wire icb_out_noearly_nxt;
  generate 
  if(WR_EARLY_RETURN == 1) begin:gen_wr_early_return_flg
  assign icb_noearly_vld_set = i_icb_cmd_valid & i_icb_cmd_ready & (i_icb_cmd_read | i_icb_cmd_attri[1]) & bus_clk_en;
  assign icb_out_noearly_nxt = i_icb_cmd_read | (i_icb_cmd_attri[1]);
  end
  else begin:gen_no_wr_early_return_flg
  assign icb_noearly_vld_set = i_icb_cmd_valid & i_icb_cmd_ready & bus_clk_en;
  assign icb_out_noearly_nxt = 1'b1;
  end
  endgenerate
  wire icb_noearly_vld_clr = i_icb_rsp_valid & i_icb_rsp_ready & icb_noearly_vld_r & bus_clk_en;
  wire icb_noearly_vld_ena = icb_noearly_vld_set | icb_noearly_vld_clr;
  wire icb_noearly_vld_nxt = icb_noearly_vld_set | (~icb_noearly_vld_clr);
e603_subsys_gnrl_dfflr #(1) icb_noearly_vld_dfflr (icb_noearly_vld_ena, icb_noearly_vld_nxt, icb_noearly_vld_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_out_flag_r;
  wire outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready & bus_clk_en;
  wire outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & bus_clk_en;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_out_flag_r = (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
  wire outs_cnt_eq0 = (outs_cnt_r == {{OUTS_CNT_W-1{1'b0}},1'b0});
  wire outs_cnt_eq1 = (outs_cnt_r == {{OUTS_CNT_W-1{1'b0}},1'b1});
  assign outs_cnt_max = (outs_cnt_r == {OUTS_CNT_W{1'b1}});
  assign i_icb_rsp_valid     = (~outs_cnt_eq0) & i_icb_rsp_valid_raw;
  assign i_icb_rsp_ready_raw = (~outs_cnt_eq0) & i_icb_rsp_ready;
  wire icb_out_noearly_r;
  wire icb_out_noearly_ena = i_icb_cmd_valid & i_icb_cmd_ready & bus_clk_en;
e603_subsys_gnrl_dfflr #(1) icb_out_noearly_dfflr (icb_out_noearly_ena, icb_out_noearly_nxt, icb_out_noearly_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire ahbl_hsel_trans_rd = (ahbl_hsel_trans & (~ahbl_hwrite));
  wire hready_out_condi;
  assign i_icb_cmd_valid = (
                 (ahbl_hsel_trans_rd & hready_out_condi & ahbl_hready_real)
               | (icb_wr_vld_r & (
                     (icb_out_flag_r & icb_out_noearly_r) ? (hready_out_condi & ahbl_hready_real) : 1'b1
                                 ) 
                 )
               ) 
               ;
  assign icb_cmd_sel = ahbl_hsel_trans | icb_wr_vld_r | ahbl_hsel_trans_busy | cmd_bypbuf_fifo_o_vld;
  assign rd_hresp_1st_err = (i_icb_rsp_err & icb_out_noearly_r) ? (~rd_hresp_1st_err_r) : 1'b0;
  wire   wait_wr_finish = (icb_out_flag_r & (~icb_out_noearly_r));
  generate 
if(WR_EARLY_RETURN == 1) begin:gen_wr_early_return
  assign hready_out_condi =
                (icb_out_flag_r ? ( 
                                icb_out_noearly_r ? (outs_cnt_eq1 & i_icb_rsp_valid) : 
                                (ahbl_hwrite & (~ahbl_hexcl_tie) & (~ahbl_hwrite_device)) ? (~outs_cnt_max) : 
                                        (outs_cnt_eq1 & i_icb_rsp_valid) 
                                 ) : 1'b1
                ) & 
                ((wait_wr_finish & (~ahbl_hwrite)) ? i_icb_rsp_valid : 1'b1) & 
                ((wait_wr_finish & ahbl_hwrite & (ahbl_hexcl_tie | ahbl_hwrite_device)) ? i_icb_rsp_valid : 1'b1) & 
                (
                  (~ahbl_hvalid_r) ? 1'b1 :
                  icb_noearly_vld_r ? (~rd_hresp_1st_err) :
                  icb_wr_vld_r ? (ahbl_hwrite & (~ahbl_hexcl_tie) & (~ahbl_hwrite_device) & (~ahbl_hwrite_device_r)) :
                  1'b1);
end
else begin:gen_no_wr_early_return
  assign hready_out_condi =
                (icb_out_flag_r ? ( 
                                icb_out_noearly_r ? (outs_cnt_eq1 & i_icb_rsp_valid) : 
                                        (outs_cnt_eq1 & i_icb_rsp_valid) 
                                 ) : 1'b1
                ) & 
                (wait_wr_finish ? i_icb_rsp_valid : 1'b1) & 
                (
                  (~ahbl_hvalid_r) ? 1'b1 :
                  icb_noearly_vld_r ? (~rd_hresp_1st_err) :
                  icb_wr_vld_r ? 1'b0 :
                  1'b1);
end
  endgenerate
  assign ahbl_hready_out = (ahbl_htrans_r == 2'b01) ? 1'b1 : (i_icb_cmd_ready & hready_out_condi); 
  assign i_icb_rsp_ready = (ahbl_hready_real & (~rd_hresp_1st_err))
                         | wait_wr_finish;
  assign ahbl_hrdata = i_icb_rsp_rdata;
  assign ahbl_hruser = i_icb_rsp_usr;
  assign ahbl_hresp[0]  = icb_noearly_vld_r ? (i_icb_rsp_err & i_icb_rsp_valid) : 1'b0;
  assign ahbl_hresp[1]  = 1'b0;
  assign ahbl_hresp_exok  = i_icb_rsp_excl_ok;
  assign ahbl2icb_active = i_icb_cmd_valid | icb_cmd_valid | icb_out_flag_r | ahbl_htrans[1];
endmodule
module e603_subsys_gnrl_ficb_active # (
  parameter OUTS_CNT_W = 1
) (
  output             icb_active,
  input              icb_cmd_valid,
  input              icb_cmd_ready,
  input              icb_rsp_valid,
  input              icb_rsp_ready,
  input              clk,
  input              rst_n
  );
  wire outs_cnt_inc = icb_cmd_valid & icb_cmd_ready
                    ;
  wire outs_cnt_dec = icb_rsp_valid & icb_rsp_ready
                    ;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_active = (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
endmodule
module e603_subsys_gnrl_usr_ficb2apb # (
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
  parameter AW = 32,
  parameter DW = 32 
) (
  input              icb_cmd_sel ,
  input              icb_cmd_valid,
  output             icb_cmd_ready,
  input              icb_cmd_read,
  input  [AW-1:0]    icb_cmd_addr,
  input  [DW-1:0]    icb_cmd_wdata,
  input  [(DW/8-1):0]  icb_cmd_wmask,
  input  [1:0]       icb_cmd_beat,
  input  [2:0]       icb_cmd_size,
  input              icb_cmd_excl,
  input              icb_cmd_lock,
  input  [7:0]       icb_cmd_xlen,
  input  [1:0]       icb_cmd_xburst,
  input  [1:0]       icb_cmd_modes,
  input              icb_cmd_dmode,
  input  [2:0]       icb_cmd_attri,
  output             icb_rsp_valid,
  input              icb_rsp_ready,
  output             icb_rsp_err,
  output             icb_rsp_excl_ok,
  output [DW-1:0]    icb_rsp_rdata,
  output [AW-1:0] apb_paddr,
  output          apb_pwrite,
  output          apb_psel,
  output [2:0]    apb_pprot,
  output [(DW/8-1):0]    apb_pstrobe,
  output          apb_penable,
  output [DW-1:0] apb_pwdata,
  input  [DW-1:0] apb_prdata,
  input           apb_pready,
  input           apb_pslverr,
  input  [CMD_UW-1:0]    icb_cmd_usr,
  output [RSP_UW-1:0]    icb_rsp_usr,
  output [CMD_UW-1:0]    apb_puser,
  input  [RSP_UW-1:0]    apb_pruser,
  input           bus_clk_en,
  input  clk,
  input  rst_n
  );
  wire            i_icb_rsp_valid;
  wire            i_icb_rsp_ready;
  wire            i_icb_rsp_err  ;
  wire            i_icb_rsp_excl_ok  ;
  wire [DW-1:0]   i_icb_rsp_rdata;
  wire [RSP_UW-1:0] i_icb_rsp_usr;
  localparam RSP_PACK_W = (2+DW
                          +RSP_UW
                     );
 wire burst_valid_r;
  wire apb_enable_r;
 wire icb_cmd_hsked = icb_cmd_valid & icb_cmd_ready;
 wire icb_cmd_ready_pre;
 wire apb_enable_set;
 wire apb_enable_clr;
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 i_icb_rsp_err,
                                 i_icb_rsp_excl_ok,
                                 i_icb_rsp_rdata 
                                ,i_icb_rsp_usr
                                 };
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 icb_rsp_err,
                                 icb_rsp_excl_ok,
                                 icb_rsp_rdata 
                                ,icb_rsp_usr
                                } = rsp_fifo_o_dat;
    assign icb_rsp_valid   = i_icb_rsp_valid; 
    assign i_icb_rsp_ready = icb_rsp_ready; 
    assign rsp_fifo_o_dat = rsp_fifo_i_dat;
    assign burst_valid_r = 1'b0;
    wire burst_valid_real = 1'b0;
  assign i_icb_rsp_valid = icb_cmd_ready_pre;
  wire i_icb_rsp_fifo_avail = 1'b1;
  assign i_icb_rsp_rdata = apb_prdata;
  assign i_icb_rsp_excl_ok = 1'b0;
  assign i_icb_rsp_err = apb_pslverr;
  assign apb_enable_set = (~apb_enable_r) & ((icb_cmd_valid & i_icb_rsp_fifo_avail & (~burst_valid_r)) | burst_valid_real);
  assign icb_cmd_ready_pre = (apb_enable_r & apb_pready);
  assign icb_cmd_ready = icb_cmd_ready_pre & (~burst_valid_r) & i_icb_rsp_fifo_avail;
  assign apb_enable_clr = icb_cmd_ready_pre;
  wire apb_enable_ena = bus_clk_en & (apb_enable_set | apb_enable_clr);
  wire apb_enable_nxt = apb_enable_set & (~apb_enable_clr);
e603_subsys_gnrl_dfflr #(1) apb_enable_dfflr (apb_enable_ena, apb_enable_nxt, apb_enable_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_cmd_mmode  = (icb_cmd_modes == 2'd0);
  wire icb_cmd_hmode  = (icb_cmd_modes == 2'd1);
  wire icb_cmd_smode  = (icb_cmd_modes == 2'd2);
  wire icb_cmd_umode  = (icb_cmd_modes == 2'd3);
  wire icb_cmd_ifu    = icb_cmd_attri[0];
  wire [AW-1:0] icb_cmd_addr_r = {AW{1'b0}};
  wire icb_cmd_mmode_r = 1'b0;
  wire icb_cmd_ifu_r = 1'b0;
  wire  [CMD_UW-1:0]    icb_cmd_usr_r = {CMD_UW{1'b0}};
  assign apb_paddr  = burst_valid_r ? icb_cmd_addr_r : icb_cmd_addr;
  assign apb_pwrite = burst_valid_r ? 1'b0 : (~icb_cmd_read);
  assign apb_pprot[0] = burst_valid_r ? icb_cmd_mmode_r : icb_cmd_mmode;
  assign apb_pprot[1] = 1'b1         ;
  assign apb_pprot[2] = burst_valid_r ? icb_cmd_ifu_r : icb_cmd_ifu  ;
  assign apb_psel    = (icb_cmd_valid & i_icb_rsp_fifo_avail & (~burst_valid_r)) | burst_valid_real | apb_enable_r;
  assign apb_penable = apb_enable_r;
  assign apb_pwdata  = (burst_valid_r | icb_cmd_read) ? {DW{1'b0}} : icb_cmd_wdata;
  assign apb_pstrobe = (burst_valid_r | icb_cmd_read) ? {DW/8{1'b0}} : icb_cmd_wmask;
  assign apb_puser  = burst_valid_r ? icb_cmd_usr_r : icb_cmd_usr;
  assign i_icb_rsp_usr = apb_pruser; 
endmodule
module e603_subsys_gnrl_apb2ficb_zero # (
  parameter AW = 32,
  parameter DW = 64 
) (
  output              icb_cmd_sel,
  output              icb_cmd_valid,
  input               icb_cmd_ready,
  output              icb_cmd_read,
  output  [AW-1:0]    icb_cmd_addr,
  output  [DW-1:0]    icb_cmd_wdata,
  output  [(DW/8-1):0]  icb_cmd_wmask,
  output  [2:0]       icb_cmd_size,
  output [7:0]       icb_cmd_xlen,
  output [1:0]       icb_cmd_xburst,
  output [1:0]       icb_cmd_modes,
  output             icb_cmd_dmode,
  output [2:0]       icb_cmd_attri,
  input               icb_rsp_valid,
  input               icb_rsp_err,
  input   [DW-1:0]    icb_rsp_rdata,
  input   [AW-1:0] apb_paddr,
  input            apb_pwrite,
  input            apb_psel ,
  input            apb_penable,
  input   [DW-1:0] apb_pwdata,
  output  [DW-1:0] apb_prdata,
  output           apb_pready,
  output           apb_pslverr,
  input  clk,
  input  rst_n
  );
  assign apb_prdata  = icb_rsp_rdata;
  assign apb_pslverr = icb_rsp_err;
  assign apb_pready    = icb_cmd_ready;
  assign icb_cmd_valid = apb_psel & apb_penable;
  assign icb_cmd_sel   = icb_cmd_valid;
  assign icb_cmd_read  = ~apb_pwrite;
  assign icb_cmd_addr  = apb_paddr;
  assign icb_cmd_wdata = apb_pwdata;
  assign icb_cmd_wmask = {DW/8{1'b1}};
  assign icb_cmd_xlen   = 8'b0;
  assign icb_cmd_xburst = 2'b0;
  assign icb_cmd_modes  = 2'b0;
  assign icb_cmd_dmode  = 1'b0;
  assign icb_cmd_attri  = 3'b0;
  generate
    if(DW == 8) begin:gen_dw8
      assign icb_cmd_size = 3'b00;
    end
    if(DW == 16) begin:gen_dw16
      assign icb_cmd_size = 3'b01;
    end
    if(DW == 32) begin:gen_dw32
      assign icb_cmd_size = 3'b10;
    end
    if(DW == 64) begin:gen_dw64
      assign icb_cmd_size = 3'b11;
    end
  endgenerate
endmodule
module e603_subsys_gnrl_usr_apb2ficb # (
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
  parameter AW = 32,
  parameter DW = 64 
) (
  input bus_clk_en,
  output apb2icb_active,
  output              icb_cmd_sel,
  output              icb_cmd_valid,
  input               icb_cmd_ready,
  output              icb_cmd_read,
  output  [AW-1:0]    icb_cmd_addr,
  output  [DW-1:0]    icb_cmd_wdata,
  output  [(DW/8-1):0]  icb_cmd_wmask,
  output  [2:0]       icb_cmd_size,
  output [7:0]       icb_cmd_xlen,
  output [1:0]       icb_cmd_xburst,
  output [1:0]       icb_cmd_modes,
  output             icb_cmd_dmode,
  output [2:0]       icb_cmd_attri,
  output              icb_cmd_lock,
  output              icb_cmd_excl,
  output [1:0]        icb_cmd_beat,
  input               icb_rsp_valid,
  output              icb_rsp_ready,
  input               icb_rsp_err,
  input   [DW-1:0]    icb_rsp_rdata,
  input               icb_rsp_excl_ok,
  output  [CMD_UW-1:0]    icb_cmd_usr,
  input   [RSP_UW-1:0]    icb_rsp_usr,
  input   [CMD_UW-1:0]    apb_puser,
  output  [RSP_UW-1:0]    apb_pruser,
  input   [AW-1:0] apb_paddr,
  input            apb_pwrite,
  input            apb_psel ,
  input            apb_penable,
  input   [DW-1:0] apb_pwdata,
  output  [DW-1:0] apb_prdata,
  output           apb_pready,
  output           apb_pslverr,
  input [2:0]    apb_pprot,
  input [(DW/8-1):0]    apb_pstrobe,
  input  clk,
  input  rst_n
  );
  assign apb_prdata  = icb_rsp_rdata;
  assign apb_pslverr = icb_rsp_err;
  assign apb_pready    = icb_rsp_valid;
  wire ongoing_r;
  assign icb_cmd_valid = (apb_psel & apb_penable) & (~ongoing_r);
  assign icb_cmd_sel   = icb_cmd_valid;
  assign icb_cmd_read  = ~apb_pwrite;
  assign icb_cmd_addr  = apb_paddr;
  assign icb_cmd_wdata = apb_pwdata;
  wire icb_cmd_mmode = apb_pprot[0];
  wire icb_cmd_ifu   = apb_pprot[2];
  assign icb_cmd_modes = icb_cmd_mmode ? 2'd0 : 2'd3; 
  assign icb_cmd_wmask = icb_cmd_read ? {DW/8{1'b0}} : apb_pstrobe;
  assign icb_cmd_attri[0] = icb_cmd_ifu   ;
  assign icb_cmd_attri[1] = 1'b0;
  assign icb_cmd_attri[2] = 1'b0;
  assign icb_cmd_xlen   = 8'b0;
  assign icb_cmd_xburst = 2'b0;
  assign icb_cmd_dmode  = 1'b0;
  assign icb_cmd_lock   = 1'b0;
  assign icb_cmd_excl   = 1'b0;
  assign icb_cmd_beat   = 2'b0;
  generate
    if(DW == 8) begin:gen_dw8
      assign icb_cmd_size = 2'b00;
    end
    if(DW == 16) begin:gen_dw16
      assign icb_cmd_size = 2'b01;
    end
    if(DW == 32) begin:gen_dw32
      assign icb_cmd_size = 2'b10;
    end
    if(DW == 64) begin:gen_dw64
      assign icb_cmd_size = 2'b11;
    end
  endgenerate
  assign icb_rsp_ready = 1'b1;
  wire icb_cmd_hsked = icb_cmd_valid & icb_cmd_ready & bus_clk_en;
  wire icb_rsp_hsked = icb_rsp_valid & icb_rsp_ready & bus_clk_en;
  wire ongoing_set = icb_cmd_hsked & (~icb_rsp_hsked);
  wire ongoing_clr = icb_rsp_hsked;
  wire ongoing_ena = (ongoing_set | ongoing_clr);
  wire ongoing_nxt = (~ongoing_clr);
e603_subsys_gnrl_dfflr #(1) ongoing_dfflr (ongoing_ena, ongoing_nxt, ongoing_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign apb2icb_active = icb_cmd_valid | ongoing_r;
  assign icb_cmd_usr = apb_puser;
  assign apb_pruser  = icb_rsp_usr;
endmodule
module e603_subsys_gnrl_usr_apb2ficb_ratio #(
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter SUPPORT_RATIO = 0,
    parameter CMD_DP = 0,
    parameter RSP_DP = 0,
    parameter RSP_BYPBUF = 0,
    parameter AW = 32,
    parameter DW = 32
)(
  output apb2icb_ratio_active,
  input  icb_clk_en,
  input  ratio_apb_clk_en,
  input  [CMD_UW              -1:0] apb_puser,
  output [RSP_UW              -1:0] apb_pruser,
  output [         RSP_UW-1:0]   icb_cmd_usr,
  input  [        RSP_UW-1:0]    icb_rsp_usr,
  input   [AW-1:0] apb_paddr,
  input            apb_pwrite,
  input            apb_psel ,
  input            apb_penable,
  input   [DW-1:0] apb_pwdata,
  output  [DW-1:0] apb_prdata,
  output           apb_pready,
  output           apb_pslverr,
  input [2:0]    apb_pprot,
  input [3:0]    apb_pstrobe,
  output                         icb_cmd_valid,
  input                          icb_cmd_ready,
  output [             AW-1:0]   icb_cmd_addr,
  output                         icb_cmd_read,
  output [        DW-1:0]        icb_cmd_wdata,
  output [        DW/8-1:0]      icb_cmd_wmask,
  output                         icb_cmd_lock,
  output                         icb_cmd_excl,
  output [2:0]                   icb_cmd_size,
  output                         icb_cmd_sel,
  output [1:0]                   icb_cmd_beat,
  output [7:0]                   icb_cmd_xlen,
  output [1:0]                   icb_cmd_xburst,
  output [1:0]                   icb_cmd_modes,
  output                         icb_cmd_dmode,
  output [2:0]                   icb_cmd_attri,
  input                          icb_rsp_valid,
  output                         icb_rsp_ready,
  input                          icb_rsp_err  ,
  input                          icb_rsp_excl_ok,
  input  [        DW-1:0]        icb_rsp_rdata,
  input  clk,
  input  rst_n
  );
  wire apb2icb_active;
  wire            buf_icb_cmd_valid;
  wire            buf_icb_cmd_ready;
  wire [AW-1:0]   buf_icb_cmd_addr;
  wire            buf_icb_cmd_read;
  wire  [1:0]     buf_icb_cmd_beat;
  wire  [7:0]     buf_icb_cmd_xlen;
  wire  [1:0]     buf_icb_cmd_xburst;
  wire  [1:0]     buf_icb_cmd_modes;
  wire            buf_icb_cmd_dmode;
  wire  [2:0]     buf_icb_cmd_attri;
  wire [DW-1:0]   buf_icb_cmd_wdata;
  wire [DW/8-1:0] buf_icb_cmd_wmask;
  wire            buf_icb_cmd_lock;
  wire            buf_icb_cmd_excl;
  wire [2:0]      buf_icb_cmd_size;
  wire            buf_icb_rsp_valid;
  wire            buf_icb_rsp_ready;
  wire            buf_icb_rsp_err  ;
  wire            buf_icb_rsp_excl_ok  ;
  wire [DW-1:0]   buf_icb_rsp_rdata;
  wire [CMD_UW-1:0]   buf_icb_cmd_usr;
  wire [RSP_UW-1:0]   buf_icb_rsp_usr;
  e603_subsys_gnrl_usr_apb2ficb
  #(
      .CMD_UW(CMD_UW),
      .RSP_UW(RSP_UW),
      .AW(AW),
      .DW(DW)
    ) u_apb2icb(
    .bus_clk_en        (ratio_apb_clk_en),
    .apb2icb_active   (apb2icb_active),
    .icb_cmd_sel       (),
    .icb_cmd_valid     (buf_icb_cmd_valid),
    .icb_cmd_ready     (buf_icb_cmd_ready),
    .icb_cmd_read      (buf_icb_cmd_read ),
    .icb_cmd_addr      (buf_icb_cmd_addr ),
    .icb_cmd_wdata     (buf_icb_cmd_wdata),
    .icb_cmd_wmask     (buf_icb_cmd_wmask),
    .icb_cmd_size      (buf_icb_cmd_size ),
    .icb_cmd_lock      (buf_icb_cmd_lock ),
    .icb_cmd_excl      (buf_icb_cmd_excl),
    .icb_cmd_beat      (buf_icb_cmd_beat  ),
    .icb_cmd_xlen      (buf_icb_cmd_xlen  ),
    .icb_cmd_xburst    (buf_icb_cmd_xburst),
    .icb_cmd_modes     (buf_icb_cmd_modes ),
    .icb_cmd_dmode     (buf_icb_cmd_dmode ),
    .icb_cmd_attri     (buf_icb_cmd_attri ),
    .icb_rsp_valid     (buf_icb_rsp_valid),
    .icb_rsp_ready     (buf_icb_rsp_ready),
    .icb_rsp_err       (buf_icb_rsp_err  ),
    .icb_rsp_rdata     (buf_icb_rsp_rdata),
    .icb_rsp_excl_ok   (buf_icb_rsp_excl_ok),
    .icb_cmd_usr       (buf_icb_cmd_usr),
    .icb_rsp_usr       (buf_icb_rsp_usr),
        .apb_puser      (apb_puser),
        .apb_pruser      (apb_pruser),
    .apb_paddr   (apb_paddr  ),
    .apb_pwrite  (apb_pwrite ),
    .apb_psel    (apb_psel   ),
    .apb_penable (apb_penable),
    .apb_pwdata  (apb_pwdata ),
    .apb_prdata  (apb_prdata ),
    .apb_pready  (apb_pready ),
    .apb_pslverr (apb_pslverr),
    .apb_pprot   (apb_pprot  ),
    .apb_pstrobe (apb_pstrobe),
    .clk         (clk  ),
    .rst_n       (rst_n)
  );
  wire buffer_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(SUPPORT_RATIO),
    .O_SUPPORT_RATIO(SUPPORT_RATIO),
    .OUTS_CNT_W   (2),
    .AW    (AW),
    .DW    (DW),
    .CMD_DP(CMD_DP),
    .RSP_DP(RSP_DP),
    .RSP_BYPBUF(RSP_BYPBUF),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(0),
    .CMD_UW (CMD_UW),
    .RSP_UW (RSP_UW)
  )u_icb_buffer(
    .i_clk_en (ratio_apb_clk_en),
    .o_clk_en (icb_clk_en),
    .icb_buffer_active      (buffer_active),
    .i_icb_cmd_sel          (buf_icb_cmd_valid),
    .i_icb_cmd_valid        (buf_icb_cmd_valid),
    .i_icb_cmd_ready        (buf_icb_cmd_ready),
    .i_icb_cmd_read         (buf_icb_cmd_read ),
    .i_icb_cmd_addr         (buf_icb_cmd_addr ),
    .i_icb_cmd_wdata        (buf_icb_cmd_wdata),
    .i_icb_cmd_wmask        (buf_icb_cmd_wmask),
    .i_icb_cmd_lock         (buf_icb_cmd_lock ),
    .i_icb_cmd_excl         (buf_icb_cmd_excl ),
    .i_icb_cmd_size         (buf_icb_cmd_size ),
    .i_icb_cmd_beat         (buf_icb_cmd_beat  ),
    .i_icb_cmd_xlen         (buf_icb_cmd_xlen  ),
    .i_icb_cmd_xburst       (buf_icb_cmd_xburst),
    .i_icb_cmd_modes        (buf_icb_cmd_modes ),
    .i_icb_cmd_dmode        (buf_icb_cmd_dmode ),
    .i_icb_cmd_attri        (buf_icb_cmd_attri ),
    .i_icb_rsp_valid        (buf_icb_rsp_valid),
    .i_icb_rsp_ready        (buf_icb_rsp_ready),
    .i_icb_rsp_err          (buf_icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (buf_icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (buf_icb_rsp_rdata),
    .o_icb_cmd_sel          (icb_cmd_sel  ),
    .o_icb_cmd_valid        (icb_cmd_valid),
    .o_icb_cmd_ready        (icb_cmd_ready),
    .o_icb_cmd_read         (icb_cmd_read ),
    .o_icb_cmd_addr         (icb_cmd_addr ),
    .o_icb_cmd_wdata        (icb_cmd_wdata),
    .o_icb_cmd_wmask        (icb_cmd_wmask),
    .o_icb_cmd_lock         (icb_cmd_lock ),
    .o_icb_cmd_size         (icb_cmd_size ),
    .o_icb_cmd_beat         (icb_cmd_beat  ),
    .o_icb_cmd_excl         (icb_cmd_excl  ),
    .o_icb_cmd_xlen         (icb_cmd_xlen  ),
    .o_icb_cmd_xburst       (icb_cmd_xburst),
    .o_icb_cmd_modes        (icb_cmd_modes ),
    .o_icb_cmd_dmode        (icb_cmd_dmode ),
    .o_icb_cmd_attri        (icb_cmd_attri ),
    .o_icb_rsp_valid        (icb_rsp_valid),
    .o_icb_rsp_ready        (icb_rsp_ready),
    .o_icb_rsp_err          (icb_rsp_err  ),
    .o_icb_rsp_rdata        (icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (icb_rsp_excl_ok),
    .i_icb_cmd_usr          (buf_icb_cmd_usr),
    .i_icb_rsp_usr          (buf_icb_rsp_usr),
    .o_icb_cmd_usr          (icb_cmd_usr),
    .o_icb_rsp_usr          (icb_rsp_usr  ),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
  assign apb2icb_ratio_active = apb2icb_active | buffer_active;
endmodule
module e603_subsys_gnrl_usr_apb2ficb_async # (
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
  parameter SYNC_DP = 2,
  parameter AW = 32,
  parameter DW = 32
)(
  output apb2icb_async_apb_active,
  output apb2icb_async_icb_active,
  input  icb_clk,
  input  icb_rst_n,
  input  async_apb_clk,
  input  async_apb_rst_n,
  input   [AW-1:0] apb_paddr,
  input            apb_pwrite,
  input            apb_psel ,
  input            apb_penable,
  input   [DW-1:0] apb_pwdata,
  output  [DW-1:0] apb_prdata,
  output           apb_pready,
  output           apb_pslverr,
  input [2:0]    apb_pprot,
  input [3:0]    apb_pstrobe,
  input  [CMD_UW              -1:0] apb_puser,
  output [RSP_UW              -1:0] apb_pruser,
  output [         RSP_UW-1:0]   icb_cmd_usr,
  input  [        RSP_UW-1:0]    icb_rsp_usr,
  output                         icb_cmd_valid,
  input                          icb_cmd_ready,
  output [             AW-1:0]   icb_cmd_addr,
  output                         icb_cmd_read,
  output [        DW-1:0]        icb_cmd_wdata,
  output [        DW/8-1:0]      icb_cmd_wmask,
  output                         icb_cmd_lock,
  output                         icb_cmd_excl,
  output [2:0]                   icb_cmd_size,
  output                         icb_cmd_sel,
  output [1:0]                   icb_cmd_beat,
  output [7:0]                   icb_cmd_xlen,
  output [1:0]                   icb_cmd_xburst,
  output [1:0]                   icb_cmd_modes,
  output                         icb_cmd_dmode,
  output [2:0]                   icb_cmd_attri,
  input                          icb_rsp_valid,
  output                         icb_rsp_ready,
  input                          icb_rsp_err  ,
  input                          icb_rsp_excl_ok,
  input  [        DW-1:0]        icb_rsp_rdata
  );
  wire icb2icb_async_i_active;
  wire icb2icb_async_o_active;
  wire apb2icb_active;
  wire            async_icb_cmd_valid;
  wire            async_icb_cmd_ready;
  wire [AW-1:0]   async_icb_cmd_addr;
  wire            async_icb_cmd_read;
  wire [DW-1:0]   async_icb_cmd_wdata;
  wire [DW/8-1:0] async_icb_cmd_wmask;
  wire [2:0]      async_icb_cmd_size;
  wire            async_icb_cmd_sel;
  wire            async_icb_cmd_lock;
  wire            async_icb_cmd_excl;
  wire  [1:0]     async_icb_cmd_beat;
  wire  [7:0]     async_icb_cmd_xlen;
  wire  [1:0]     async_icb_cmd_xburst;
  wire  [1:0]     async_icb_cmd_modes;
  wire            async_icb_cmd_dmode;
  wire  [2:0]     async_icb_cmd_attri;
  wire            async_icb_rsp_valid;
  wire            async_icb_rsp_ready;
  wire            async_icb_rsp_err  ;
  wire            async_icb_rsp_excl_ok  ;
  wire [DW-1:0]   async_icb_rsp_rdata;
  wire [CMD_UW-1:0]   async_icb_cmd_usr;
  wire [RSP_UW-1:0]   async_icb_rsp_usr;
  e603_subsys_gnrl_usr_apb2ficb
  #(
      .CMD_UW(CMD_UW),
      .RSP_UW(RSP_UW),
      .AW(AW),
      .DW(DW)
    ) u_apb2icb(
    .bus_clk_en        (1'b1),
    .apb2icb_active   (apb2icb_active),
    .icb_cmd_sel       (   ),
    .icb_cmd_valid     (async_icb_cmd_valid),
    .icb_cmd_ready     (async_icb_cmd_ready),
    .icb_cmd_read      (async_icb_cmd_read ),
    .icb_cmd_addr      (async_icb_cmd_addr ),
    .icb_cmd_wdata     (async_icb_cmd_wdata),
    .icb_cmd_wmask     (async_icb_cmd_wmask),
    .icb_cmd_size      (async_icb_cmd_size ),
    .icb_cmd_lock      (async_icb_cmd_lock ),
    .icb_cmd_excl      (async_icb_cmd_excl),
    .icb_cmd_beat      (async_icb_cmd_beat  ),
    .icb_cmd_xlen      (async_icb_cmd_xlen  ),
    .icb_cmd_xburst    (async_icb_cmd_xburst),
    .icb_cmd_modes     (async_icb_cmd_modes ),
    .icb_cmd_dmode     (async_icb_cmd_dmode ),
    .icb_cmd_attri     (async_icb_cmd_attri ),
    .icb_rsp_valid     (async_icb_rsp_valid),
    .icb_rsp_ready     (async_icb_rsp_ready),
    .icb_rsp_err       (async_icb_rsp_err  ),
    .icb_rsp_rdata     (async_icb_rsp_rdata),
    .icb_rsp_excl_ok   (async_icb_rsp_excl_ok),
    .icb_cmd_usr       (async_icb_cmd_usr),
    .icb_rsp_usr       (async_icb_rsp_usr),
        .apb_puser      (apb_puser),
        .apb_pruser     (apb_pruser),
    .apb_paddr   (apb_paddr  ),
    .apb_pwrite  (apb_pwrite ),
    .apb_psel    (apb_psel   ),
    .apb_penable (apb_penable),
    .apb_pwdata  (apb_pwdata ),
    .apb_prdata  (apb_prdata ),
    .apb_pready  (apb_pready ),
    .apb_pslverr (apb_pslverr),
    .apb_pprot   (apb_pprot  ),
    .apb_pstrobe (apb_pstrobe),
    .clk               (async_apb_clk  ),
    .rst_n             (async_apb_rst_n)
  );
  e603_subsys_gnrl_ficb_async # (
    .RSP_ALWAYS_READY(0),
    .OUTS_CNT_W(2),
    .SYNC_DP (SYNC_DP),
    .ASYNC_FIFO (0),
    .ASYNC_FIFO_DP(0),
    .ASYNC_FIFO_DP_PTR_W(0),
    .AW    (AW),
    .DW    (DW),
    .CMD_UW (CMD_UW),
    .RSP_UW (RSP_UW)
  )u_icb2icb_async(
    .icb2icb_async_i_active   (icb2icb_async_i_active),
    .icb2icb_async_o_active   (icb2icb_async_o_active),
    .i_clk                  (async_apb_clk),
    .i_rst_n                (async_apb_rst_n),
    .o_clk                  (icb_clk),
    .o_rst_n                (icb_rst_n),
    .i_icb_cmd_sel          (async_icb_cmd_valid),
    .i_icb_cmd_valid        (async_icb_cmd_valid),
    .i_icb_cmd_ready        (async_icb_cmd_ready),
    .i_icb_cmd_read         (async_icb_cmd_read ),
    .i_icb_cmd_addr         (async_icb_cmd_addr ),
    .i_icb_cmd_wdata        (async_icb_cmd_wdata),
    .i_icb_cmd_wmask        (async_icb_cmd_wmask),
    .i_icb_cmd_lock         (async_icb_cmd_lock   ),
    .i_icb_cmd_excl         (async_icb_cmd_excl   ),
    .i_icb_cmd_size         (async_icb_cmd_size   ),
    .i_icb_cmd_beat         (async_icb_cmd_beat   ),
    .i_icb_cmd_xlen         (async_icb_cmd_xlen   ),
    .i_icb_cmd_xburst       (async_icb_cmd_xburst ),
    .i_icb_cmd_modes        (async_icb_cmd_modes ),
    .i_icb_cmd_dmode        (async_icb_cmd_dmode ),
    .i_icb_cmd_attri        (async_icb_cmd_attri ),
    .i_icb_rsp_valid        (async_icb_rsp_valid),
    .i_icb_rsp_ready        (async_icb_rsp_ready),
    .i_icb_rsp_err          (async_icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (async_icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (async_icb_rsp_rdata),
    .i_icb_cmd_usr          (async_icb_cmd_usr),
    .i_icb_rsp_usr          (async_icb_rsp_usr),
    .o_icb_cmd_usr          (icb_cmd_usr),
    .o_icb_rsp_usr          (icb_rsp_usr  ),
    .o_icb_cmd_sel       (icb_cmd_sel  ),
    .o_icb_cmd_valid     (icb_cmd_valid),
    .o_icb_cmd_ready     (icb_cmd_ready),
    .o_icb_cmd_read      (icb_cmd_read ),
    .o_icb_cmd_addr      (icb_cmd_addr ),
    .o_icb_cmd_wdata     (icb_cmd_wdata),
    .o_icb_cmd_wmask     (icb_cmd_wmask),
    .o_icb_cmd_size      (icb_cmd_size ),
    .o_icb_cmd_beat      (icb_cmd_beat  ),
    .o_icb_cmd_lock      (icb_cmd_lock  ),
    .o_icb_cmd_excl      (icb_cmd_excl  ),
    .o_icb_cmd_xlen      (icb_cmd_xlen  ),
    .o_icb_cmd_xburst    (icb_cmd_xburst),
    .o_icb_cmd_modes     (icb_cmd_modes ),
    .o_icb_cmd_dmode     (icb_cmd_dmode ),
    .o_icb_cmd_attri     (icb_cmd_attri ),
    .o_icb_rsp_valid        (icb_rsp_valid),
    .o_icb_rsp_ready        (icb_rsp_ready),
    .o_icb_rsp_err          (icb_rsp_err  ),
    .o_icb_rsp_rdata        (icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (icb_rsp_excl_ok) 
  );
 assign apb2icb_async_apb_active = icb2icb_async_i_active | apb2icb_active;
 assign apb2icb_async_icb_active = icb2icb_async_o_active;
endmodule
module e603_subsys_gnrl_usr_ficb2apb_ratio # (
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter OUTS_CNT_W = 4,
  parameter SUPPORT_RATIO = 0,
  parameter CMD_DP = 0,
  parameter RSP_DP = 0,
  parameter RSP_BYPBUF = 0,
  parameter AW = 32,
  parameter DW = 32
)(
  output icb2apb_ratio_active,
  input  icb_clk_en,
  input  ratio_apb_clk_en,
  input              icb_cmd_excl ,
  input              icb_cmd_lock ,
  input              icb_cmd_sel ,
  input  [1:0]       icb_cmd_beat,
  input  [7:0]       icb_cmd_xlen,
  input  [1:0]       icb_cmd_xburst,
  input  [1:0]       icb_cmd_modes,
  input              icb_cmd_dmode,
  input  [2:0]       icb_cmd_attri,
  input                          icb_cmd_valid,
  output                         icb_cmd_ready,
  input  [             AW-1:0]   icb_cmd_addr,
  input                          icb_cmd_read,
  input  [        DW-1:0]        icb_cmd_wdata,
  input  [        DW/8-1:0]      icb_cmd_wmask,
  input  [2:0]                   icb_cmd_size,
  output                         icb_rsp_valid,
  input                          icb_rsp_ready,
  output                         icb_rsp_err  ,
  output                         icb_rsp_excl_ok,
  output [        DW-1:0]        icb_rsp_rdata,
  output [AW-1:0] ratio_apb_paddr,
  output          ratio_apb_pwrite,
  output          ratio_apb_psel,
  output [2:0]    ratio_apb_pprot,
  output [3:0]    ratio_apb_pstrobe,
  output          ratio_apb_penable,
  output [DW-1:0] ratio_apb_pwdata,
  input  [DW-1:0] ratio_apb_prdata,
  input           ratio_apb_pready,
  input           ratio_apb_pslverr,
  input  [CMD_UW -1:0] icb_cmd_usr,
  output [RSP_UW -1:0] icb_rsp_usr,
  output [CMD_UW              -1:0] ratio_apb_puser,
  input  [RSP_UW              -1:0] ratio_apb_pruser,
  input  clk,
  input  rst_n
  );
  wire buffer_active;
  assign icb2apb_ratio_active = buffer_active;
  wire            buf_icb_cmd_sel ;
  wire  [1:0]     buf_icb_cmd_modes;
  wire            buf_icb_cmd_dmode;
  wire  [2:0]     buf_icb_cmd_attri;
  wire            buf_icb_cmd_valid;
  wire            buf_icb_cmd_ready;
  wire [AW-1:0]   buf_icb_cmd_addr;
  wire            buf_icb_cmd_read;
  wire [DW-1:0]   buf_icb_cmd_wdata;
  wire [DW/8-1:0] buf_icb_cmd_wmask;
  wire            buf_icb_cmd_lock;
  wire            buf_icb_cmd_excl;
  wire  [1:0]     buf_icb_cmd_beat;
  wire  [7:0]     buf_icb_cmd_xlen;
  wire  [1:0]     buf_icb_cmd_xburst;
  wire [2:0]      buf_icb_cmd_size;
  wire            buf_icb_rsp_valid;
  wire            buf_icb_rsp_ready;
  wire            buf_icb_rsp_err  ;
  wire            buf_icb_rsp_excl_ok  ;
  wire [DW-1:0]   buf_icb_rsp_rdata;
  wire [CMD_UW-1:0]   buf_icb_cmd_usr;
  wire [RSP_UW-1:0]   buf_icb_rsp_usr;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(SUPPORT_RATIO),
    .O_SUPPORT_RATIO(SUPPORT_RATIO),
    .OUTS_CNT_W   (OUTS_CNT_W),
    .AW    (AW),
    .DW    (DW),
    .CMD_DP(CMD_DP),
    .RSP_DP(RSP_DP),
    .RSP_BYPBUF(RSP_BYPBUF),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(1),
    .CMD_UW (CMD_UW
            ),
    .RSP_UW (RSP_UW)
  )u_icb_buffer(
    .i_clk_en (icb_clk_en),
    .o_clk_en (ratio_apb_clk_en),
    .icb_buffer_active      (buffer_active),
    .i_icb_cmd_sel          (icb_cmd_valid),
    .i_icb_cmd_valid        (icb_cmd_valid),
    .i_icb_cmd_ready        (icb_cmd_ready),
    .i_icb_cmd_read         (icb_cmd_read ),
    .i_icb_cmd_addr         (icb_cmd_addr ),
    .i_icb_cmd_wdata        (icb_cmd_wdata),
    .i_icb_cmd_wmask        (icb_cmd_wmask),
    .i_icb_cmd_lock         (icb_cmd_lock),
    .i_icb_cmd_excl         (icb_cmd_excl),
    .i_icb_cmd_size         (icb_cmd_size ),
    .i_icb_cmd_beat         (icb_cmd_beat ),
    .i_icb_cmd_xlen         (icb_cmd_xlen    ),
    .i_icb_cmd_xburst       (icb_cmd_xburst),
    .i_icb_cmd_modes        (icb_cmd_modes  ),
    .i_icb_cmd_dmode        (icb_cmd_dmode  ),
    .i_icb_cmd_attri        (icb_cmd_attri  ),
    .i_icb_rsp_valid        (icb_rsp_valid),
    .i_icb_rsp_ready        (icb_rsp_ready),
    .i_icb_rsp_err          (icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (icb_rsp_rdata),
    .i_icb_cmd_usr          ({icb_cmd_usr
                             }
                            ),
    .i_icb_rsp_usr          (icb_rsp_usr),
    .o_icb_cmd_usr          ({buf_icb_cmd_usr
                             }
                            ),
    .o_icb_rsp_usr          (buf_icb_rsp_usr),
    .o_icb_cmd_sel          (),
    .o_icb_cmd_valid        (buf_icb_cmd_valid),
    .o_icb_cmd_ready        (buf_icb_cmd_ready),
    .o_icb_cmd_read         (buf_icb_cmd_read ),
    .o_icb_cmd_addr         (buf_icb_cmd_addr ),
    .o_icb_cmd_wdata        (buf_icb_cmd_wdata),
    .o_icb_cmd_wmask        (buf_icb_cmd_wmask),
    .o_icb_cmd_lock         (buf_icb_cmd_lock ),
    .o_icb_cmd_size         (buf_icb_cmd_size ),
    .o_icb_cmd_beat         (buf_icb_cmd_beat  ),
    .o_icb_cmd_excl         (buf_icb_cmd_excl  ),
    .o_icb_cmd_xlen         (buf_icb_cmd_xlen    ),
    .o_icb_cmd_xburst       (buf_icb_cmd_xburst),
    .o_icb_cmd_modes        (buf_icb_cmd_modes ),
    .o_icb_cmd_dmode        (buf_icb_cmd_dmode ),
    .o_icb_cmd_attri        (buf_icb_cmd_attri ),
    .o_icb_rsp_valid        (buf_icb_rsp_valid),
    .o_icb_rsp_ready        (buf_icb_rsp_ready),
    .o_icb_rsp_err          (buf_icb_rsp_err  ),
    .o_icb_rsp_rdata        (buf_icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (buf_icb_rsp_excl_ok),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
  e603_subsys_gnrl_usr_ficb2apb
  #(
      .CMD_UW(CMD_UW),
    .RSP_UW(RSP_UW),
  .AW(AW),
  .DW(DW)
  ) u_e603_subsys_gnrl_ficb2apb(
    .icb_cmd_sel   (buf_icb_cmd_valid ),
    .icb_cmd_valid (buf_icb_cmd_valid ),
    .icb_cmd_ready (buf_icb_cmd_ready ),
    .icb_cmd_read  (buf_icb_cmd_read  ),
    .icb_cmd_addr  (buf_icb_cmd_addr  ),
    .icb_cmd_wdata (buf_icb_cmd_wdata ),
    .icb_cmd_wmask (buf_icb_cmd_wmask ),
    .icb_cmd_size  (buf_icb_cmd_size  ),
    .icb_cmd_excl  (buf_icb_cmd_excl   ),
    .icb_cmd_lock  (buf_icb_cmd_lock   ),
    .icb_cmd_beat  (buf_icb_cmd_beat   ),
    .icb_cmd_xlen  (buf_icb_cmd_xlen   ),
    .icb_cmd_xburst(buf_icb_cmd_xburst),
    .icb_cmd_modes (buf_icb_cmd_modes ),
    .icb_cmd_dmode (buf_icb_cmd_dmode ),
    .icb_cmd_attri (buf_icb_cmd_attri ),
    .icb_rsp_valid (buf_icb_rsp_valid ),
    .icb_rsp_err   (buf_icb_rsp_err   ),
    .icb_rsp_ready  (buf_icb_rsp_ready   ),
    .icb_rsp_excl_ok(buf_icb_rsp_excl_ok),
    .icb_rsp_rdata (buf_icb_rsp_rdata ),
    .apb_paddr     (ratio_apb_paddr     ),
    .apb_pwrite    (ratio_apb_pwrite    ),
    .apb_psel      (ratio_apb_psel      ),
    .apb_pprot     (ratio_apb_pprot     ),
    .apb_pstrobe   (ratio_apb_pstrobe   ),
    .apb_penable   (ratio_apb_penable   ),
    .apb_pwdata    (ratio_apb_pwdata    ),
    .apb_prdata    (ratio_apb_prdata    ),
    .apb_pready    (ratio_apb_pready    ),
    .apb_pslverr   (ratio_apb_pslverr   ),
    .icb_cmd_usr      (buf_icb_cmd_usr ),
    .icb_rsp_usr      (buf_icb_rsp_usr ),
    .apb_puser        (ratio_apb_puser   ),
    .apb_pruser       (ratio_apb_pruser   ),
    .bus_clk_en    (ratio_apb_clk_en    ),
    .clk   (clk  ),
    .rst_n (rst_n)
  );
endmodule
module e603_subsys_gnrl_usr_ficb2apb_async # (
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter OUTS_CNT_W = 4,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 1,
  parameter ASYNC_FIFO_DP = 4,
  parameter ASYNC_FIFO_DP_PTR_W = 2,
  parameter AW = 32,
  parameter DW = 32
)(
  output icb2apb_async_icb_active,
  output icb2apb_async_apb_active,
  input  icb_clk,
  input  icb_rst_n,
  input  async_apb_clk,
  input  async_apb_rst_n,
  input              icb_cmd_excl ,
  input              icb_cmd_lock ,
  input              icb_cmd_sel ,
  input  [1:0]       icb_cmd_beat,
  input  [7:0]       icb_cmd_xlen,
  input  [1:0]       icb_cmd_xburst,
  input  [1:0]       icb_cmd_modes,
  input              icb_cmd_dmode,
  input  [2:0]       icb_cmd_attri,
  input             icb_cmd_valid,
  output            icb_cmd_ready,
  input  [AW-1:0]   icb_cmd_addr,
  input             icb_cmd_read,
  input  [DW-1:0]   icb_cmd_wdata,
  input  [DW/8-1:0] icb_cmd_wmask,
  input  [2:0]      icb_cmd_size,
  output            icb_rsp_valid,
  input             icb_rsp_ready,
  output            icb_rsp_err,
  output            icb_rsp_excl_ok,
  output [DW-1:0]   icb_rsp_rdata,
  input  [CMD_UW -1:0] icb_cmd_usr,
  output [RSP_UW -1:0] icb_rsp_usr,
  output [CMD_UW              -1:0] async_apb_puser,
  input  [RSP_UW              -1:0] async_apb_pruser,
  output [AW-1:0] async_apb_paddr,
  output          async_apb_pwrite,
  output          async_apb_psel,
  output [2:0]    async_apb_pprot,
  output [3:0]    async_apb_pstrobe,
  output          async_apb_penable,
  output [DW-1:0] async_apb_pwdata,
  input  [DW-1:0] async_apb_prdata,
  input           async_apb_pready,
  input           async_apb_pslverr
  );
  wire icb2icb_async_i_active;
  wire icb2icb_async_o_active;
  wire            async_icb_cmd_sel ;
  wire  [1:0]     async_icb_cmd_modes;
  wire            async_icb_cmd_dmode;
  wire  [2:0]     async_icb_cmd_attri;
  wire            async_icb_cmd_valid;
  wire            async_icb_cmd_ready;
  wire [AW-1:0]   async_icb_cmd_addr;
  wire            async_icb_cmd_read;
  wire [DW-1:0]   async_icb_cmd_wdata;
  wire [DW/8-1:0] async_icb_cmd_wmask;
  wire [2:0]      async_icb_cmd_size;
  wire            async_icb_cmd_lock;
  wire            async_icb_cmd_excl;
  wire  [1:0]     async_icb_cmd_beat;
  wire  [7:0]     async_icb_cmd_xlen;
  wire  [1:0]     async_icb_cmd_xburst;
  wire            async_icb_rsp_valid;
  wire            async_icb_rsp_ready;
  wire            async_icb_rsp_err  ;
  wire            async_icb_rsp_excl_ok  ;
  wire [DW-1:0]   async_icb_rsp_rdata;
  wire [CMD_UW-1:0]   async_icb_cmd_usr;
  wire [RSP_UW-1:0]   async_icb_rsp_usr;
  wire [CMD_UW-1:0]   o_icb_cmd_usr;
  wire [RSP_UW-1:0]   o_icb_rsp_usr;
  wire            o_icb_cmd_sel ;
  wire  [1:0]     o_icb_cmd_modes;
  wire            o_icb_cmd_dmode;
  wire  [2:0]     o_icb_cmd_attri;
  wire            o_icb_cmd_valid;
  wire            o_icb_cmd_ready;
  wire [AW-1:0]   o_icb_cmd_addr;
  wire            o_icb_cmd_read;
  wire [DW-1:0]   o_icb_cmd_wdata;
  wire [DW/8-1:0] o_icb_cmd_wmask;
  wire [2:0]      o_icb_cmd_size;
  wire            o_icb_cmd_lock;
  wire            o_icb_cmd_excl;
  wire  [1:0]     o_icb_cmd_beat;
  wire  [7:0]     o_icb_cmd_xlen;
  wire  [1:0]     o_icb_cmd_xburst;
  wire            o_icb_rsp_valid;
  wire            o_icb_rsp_ready;
  wire            o_icb_rsp_err  ;
  wire            o_icb_rsp_excl_ok  ;
  wire [DW-1:0]   o_icb_rsp_rdata;
  e603_subsys_gnrl_ficb_async # (
    .RSP_ALWAYS_READY(0),
    .OUTS_CNT_W(OUTS_CNT_W),
    .SYNC_DP (SYNC_DP),
    .ASYNC_FIFO   (ASYNC_FIFO   ),
    .ASYNC_FIFO_DP(ASYNC_FIFO_DP),
    .ASYNC_FIFO_DP_PTR_W(ASYNC_FIFO_DP_PTR_W),
    .AW    (AW),
    .DW    (DW),
    .CMD_UW (CMD_UW
            ),
    .RSP_UW (RSP_UW)
  )u_icb2icb_async(
    .icb2icb_async_i_active   (icb2icb_async_i_active),
    .icb2icb_async_o_active   (icb2icb_async_o_active),
    .i_clk                  (icb_clk),
    .i_rst_n                (icb_rst_n),
    .i_icb_cmd_sel          (icb_cmd_valid),
    .i_icb_cmd_valid        (icb_cmd_valid),
    .i_icb_cmd_ready        (icb_cmd_ready),
    .i_icb_cmd_read         (icb_cmd_read ),
    .i_icb_cmd_addr         (icb_cmd_addr ),
    .i_icb_cmd_wdata        (icb_cmd_wdata),
    .i_icb_cmd_wmask        (icb_cmd_wmask),
    .i_icb_cmd_lock         (icb_cmd_lock),
    .i_icb_cmd_excl         (icb_cmd_excl),
    .i_icb_cmd_size         (icb_cmd_size ),
    .i_icb_cmd_beat         (icb_cmd_beat),
    .i_icb_cmd_xlen         (icb_cmd_xlen    ),
    .i_icb_cmd_xburst       (icb_cmd_xburst),
    .i_icb_cmd_modes        (icb_cmd_modes  ),
    .i_icb_cmd_dmode        (icb_cmd_dmode  ),
    .i_icb_cmd_attri        (icb_cmd_attri  ),
    .i_icb_rsp_valid        (icb_rsp_valid),
    .i_icb_rsp_ready        (icb_rsp_ready),
    .i_icb_rsp_err          (icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (icb_rsp_rdata),
    .o_clk                  (async_apb_clk),
    .o_rst_n                (async_apb_rst_n),
    .i_icb_cmd_usr          ({icb_cmd_usr
                             }
                            ),
    .i_icb_rsp_usr          (icb_rsp_usr),
    .o_icb_cmd_usr          ({async_icb_cmd_usr
                             }
                            ),
    .o_icb_rsp_usr          (async_icb_rsp_usr),
    .o_icb_cmd_sel          (),
    .o_icb_cmd_valid        (async_icb_cmd_valid),
    .o_icb_cmd_ready        (async_icb_cmd_ready),
    .o_icb_cmd_read         (async_icb_cmd_read ),
    .o_icb_cmd_addr         (async_icb_cmd_addr ),
    .o_icb_cmd_wdata        (async_icb_cmd_wdata),
    .o_icb_cmd_wmask        (async_icb_cmd_wmask),
    .o_icb_cmd_lock         (async_icb_cmd_lock),
    .o_icb_cmd_size         (async_icb_cmd_size ),
    .o_icb_cmd_beat         (async_icb_cmd_beat  ),
    .o_icb_cmd_excl         (async_icb_cmd_excl  ),
    .o_icb_cmd_xlen         (async_icb_cmd_xlen  ),
    .o_icb_cmd_xburst       (async_icb_cmd_xburst),
    .o_icb_cmd_modes        (async_icb_cmd_modes ),
    .o_icb_cmd_dmode        (async_icb_cmd_dmode ),
    .o_icb_cmd_attri        (async_icb_cmd_attri ),
    .o_icb_rsp_valid        (async_icb_rsp_valid),
    .o_icb_rsp_ready        (async_icb_rsp_ready),
    .o_icb_rsp_err          (async_icb_rsp_err  ),
    .o_icb_rsp_rdata        (async_icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (async_icb_rsp_excl_ok) 
  );
  wire o_buffer_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(0),
    .O_SUPPORT_RATIO(0),
    .AW    (AW),
    .DW    (DW),
    .CMD_DP(0),
    .RSP_BYPBUF(1),
    .RSP_DP(2),
    .OUTS_CNT_W   (2),
    .RSP_ALWAYS_READY(1),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .CMD_UW (CMD_UW
            ),
    .RSP_UW (RSP_UW)
  )u_icb_buffer(
    .i_clk_en (1'b1),
    .o_clk_en (1'b1),
    .icb_buffer_active      (o_buffer_active),
    .i_icb_cmd_sel          (async_icb_cmd_valid),
    .i_icb_cmd_valid        (async_icb_cmd_valid),
    .i_icb_cmd_ready        (async_icb_cmd_ready),
    .i_icb_cmd_read         (async_icb_cmd_read ),
    .i_icb_cmd_addr         (async_icb_cmd_addr ),
    .i_icb_cmd_wdata        (async_icb_cmd_wdata),
    .i_icb_cmd_wmask        (async_icb_cmd_wmask),
    .i_icb_cmd_lock         (async_icb_cmd_lock),
    .i_icb_cmd_excl         (async_icb_cmd_excl),
    .i_icb_cmd_size         (async_icb_cmd_size ),
    .i_icb_cmd_beat         (async_icb_cmd_beat),
    .i_icb_cmd_xlen         (async_icb_cmd_xlen    ),
    .i_icb_cmd_xburst       (async_icb_cmd_xburst),
    .i_icb_cmd_modes        (async_icb_cmd_modes ),
    .i_icb_cmd_dmode        (async_icb_cmd_dmode ),
    .i_icb_cmd_attri        (async_icb_cmd_attri ),
    .i_icb_rsp_valid        (async_icb_rsp_valid),
    .i_icb_rsp_ready        (async_icb_rsp_ready),
    .i_icb_rsp_err          (async_icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (async_icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (async_icb_rsp_rdata),
    .i_icb_cmd_usr          ({async_icb_cmd_usr
                             }
                            ),
    .i_icb_rsp_usr          (async_icb_rsp_usr),
    .o_icb_cmd_usr          ({o_icb_cmd_usr
                             }
                            ),
    .o_icb_rsp_usr          (o_icb_rsp_usr),
    .o_icb_cmd_sel          (),
    .o_icb_cmd_valid        (o_icb_cmd_valid),
    .o_icb_cmd_ready        (o_icb_cmd_ready),
    .o_icb_cmd_read         (o_icb_cmd_read ),
    .o_icb_cmd_addr         (o_icb_cmd_addr ),
    .o_icb_cmd_wdata        (o_icb_cmd_wdata),
    .o_icb_cmd_wmask        (o_icb_cmd_wmask),
    .o_icb_cmd_lock         (o_icb_cmd_lock),
    .o_icb_cmd_size         (o_icb_cmd_size ),
    .o_icb_cmd_beat         (o_icb_cmd_beat  ),
    .o_icb_cmd_excl         (o_icb_cmd_excl  ),
    .o_icb_cmd_xlen         (o_icb_cmd_xlen  ),
    .o_icb_cmd_xburst       (o_icb_cmd_xburst),
    .o_icb_cmd_modes        (o_icb_cmd_modes ),
    .o_icb_cmd_dmode        (o_icb_cmd_dmode ),
    .o_icb_cmd_attri        (o_icb_cmd_attri ),
    .o_icb_rsp_valid        (o_icb_rsp_valid),
    .o_icb_rsp_ready        (o_icb_rsp_ready),
    .o_icb_rsp_err          (o_icb_rsp_err  ),
    .o_icb_rsp_rdata        (o_icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (o_icb_rsp_excl_ok),
    .clk   (async_apb_clk  ),
    .rst_n (async_apb_rst_n)
  );
  e603_subsys_gnrl_usr_ficb2apb
  #(
    .CMD_UW(CMD_UW),
    .RSP_UW(RSP_UW),
  .AW(AW),
  .DW(DW)
  ) u_e603_subsys_gnrl_ficb2apb(
    .icb_cmd_sel   (o_icb_cmd_valid ),
    .icb_cmd_valid (o_icb_cmd_valid ),
    .icb_cmd_ready (o_icb_cmd_ready ),
    .icb_cmd_read  (o_icb_cmd_read  ),
    .icb_cmd_addr  (o_icb_cmd_addr  ),
    .icb_cmd_wdata (o_icb_cmd_wdata ),
    .icb_cmd_wmask (o_icb_cmd_wmask ),
    .icb_cmd_size  (o_icb_cmd_size  ),
    .icb_cmd_xlen  (o_icb_cmd_xlen  ),
    .icb_cmd_excl  (o_icb_cmd_excl  ),
    .icb_cmd_lock  (o_icb_cmd_lock  ),
    .icb_cmd_beat  (o_icb_cmd_beat  ),
    .icb_cmd_xburst(o_icb_cmd_xburst),
    .icb_cmd_modes (o_icb_cmd_modes ),
    .icb_cmd_dmode (o_icb_cmd_dmode ),
    .icb_cmd_attri (o_icb_cmd_attri ),
    .icb_rsp_valid (o_icb_rsp_valid ),
    .icb_rsp_err   (o_icb_rsp_err   ),
    .icb_rsp_ready (o_icb_rsp_ready   ),
    .icb_rsp_excl_ok (o_icb_rsp_excl_ok),
    .icb_rsp_rdata (o_icb_rsp_rdata ),
    .icb_cmd_usr      (o_icb_cmd_usr ),
    .icb_rsp_usr      (o_icb_rsp_usr ),
    .apb_puser        (async_apb_puser   ),
    .apb_pruser       (async_apb_pruser   ),
    .apb_paddr     (async_apb_paddr     ),
    .apb_pwrite    (async_apb_pwrite    ),
    .apb_psel      (async_apb_psel      ),
    .apb_pprot     (async_apb_pprot     ),
    .apb_pstrobe   (async_apb_pstrobe   ),
    .apb_penable   (async_apb_penable   ),
    .apb_pwdata    (async_apb_pwdata    ),
    .apb_prdata    (async_apb_prdata    ),
    .apb_pready    (async_apb_pready    ),
    .apb_pslverr   (async_apb_pslverr   ),
    .bus_clk_en    (1'b1    ),
    .clk   (async_apb_clk  ),
    .rst_n (async_apb_rst_n)
  );
 assign icb2apb_async_icb_active = icb2icb_async_i_active;
 assign icb2apb_async_apb_active = icb2icb_async_o_active | o_buffer_active;
endmodule
module e603_subsys_gnrl_usr_ficb2ahbl_ratio #(
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter OUTS_CNT_W = 2,
    parameter MON_DATA_WIDTH = 2,
    parameter SUPPORT_RATIO = 0,
    parameter CMD_DP = 0,
    parameter RSP_DP = 2,
    parameter RSP_BYPBUF = 1,
    parameter AW = 32,
    parameter DW = 32
)(
  output icb2ahbl_ratio_active,
  output icb2ahbl_pend_active,
  input  icb_clk_en,
  input  ratio_ahbl_clk_en,
  input  [CMD_UW -1:0] icb_cmd_usr,
  output [RSP_UW -1:0] icb_rsp_usr,
  output [CMD_UW              -1:0] ratio_huser,
  input  [RSP_UW              -1:0] ratio_hruser,
  input                          icb_cmd_valid,
  output                         icb_cmd_ready,
  input  [             AW-1:0]   icb_cmd_addr,
  input                          icb_cmd_read,
  input  [        DW-1:0]        icb_cmd_wdata,
  input  [        DW/8-1:0]      icb_cmd_wmask,
  input                          icb_cmd_lock,
  input                          icb_cmd_excl,
  input  [2:0]                   icb_cmd_size,
  input                          icb_cmd_sel,
  input  [1:0]                   icb_cmd_beat,
  input  [7:0]                   icb_cmd_xlen,
  input  [1:0]                   icb_cmd_xburst,
  input  [1:0]                   icb_cmd_modes,
  input                          icb_cmd_dmode,
  input  [2:0]                   icb_cmd_attri,
  output                         icb_rsp_valid,
  input                          icb_rsp_ready,
  output                         icb_rsp_err  ,
  output                         icb_rsp_excl_ok,
  output [        DW-1:0]        icb_rsp_rdata,
  output [1:0]                      ratio_htrans,
  output                            ratio_hwrite,
  output                            ratio_hmastlock,
  output [2:0]                      ratio_hsize,
  output [2:0]                      ratio_hburst,
  output [3:0]                      ratio_hprot,
  output [DW                  -1:0] ratio_hwdata,
  output [AW                  -1:0] ratio_haddr,
  input  [DW                  -1:0] ratio_hrdata,
  input  [1:0]                      ratio_hresp,
  input                             ratio_hready,
  input  clk,
  input  rst_n
  );
  wire buffer_active;
  wire            buf_icb_cmd_valid;
  wire            buf_icb_cmd_ready;
  wire [AW-1:0]   buf_icb_cmd_addr;
  wire            buf_icb_cmd_read;
  wire  [1:0]     buf_icb_cmd_beat;
  wire  [7:0]     buf_icb_cmd_xlen;
  wire  [1:0]     buf_icb_cmd_xburst;
  wire  [1:0]     buf_icb_cmd_modes;
  wire            buf_icb_cmd_dmode;
  wire  [2:0]     buf_icb_cmd_attri;
  wire [DW-1:0]   buf_icb_cmd_wdata;
  wire [DW/8-1:0] buf_icb_cmd_wmask;
  wire            buf_icb_cmd_lock;
  wire            buf_icb_cmd_excl;
  wire [2:0]      buf_icb_cmd_size;
  wire            buf_icb_rsp_valid;
  wire            buf_icb_rsp_ready;
  wire            buf_icb_rsp_err  ;
  wire            buf_icb_rsp_excl_ok  ;
  wire [DW-1:0]   buf_icb_rsp_rdata;
  wire [CMD_UW-1:0]   buf_icb_cmd_usr;
  wire [RSP_UW-1:0]   buf_icb_rsp_usr;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(SUPPORT_RATIO),
    .O_SUPPORT_RATIO(SUPPORT_RATIO),
    .OUTS_CNT_W   (OUTS_CNT_W),
    .AW    (AW),
    .DW    (DW),
    .CMD_DP(CMD_DP),
    .RSP_DP(RSP_DP),
    .RSP_BYPBUF(RSP_BYPBUF),
        .RSP_ALWAYS_READY(1),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .CMD_UW (CMD_UW),
    .RSP_UW (RSP_UW)
  )u_icb_buffer(
    .i_clk_en (icb_clk_en),
    .o_clk_en (ratio_ahbl_clk_en),
    .icb_buffer_active      (buffer_active),
    .i_icb_cmd_sel          (icb_cmd_valid),
    .i_icb_cmd_valid        (icb_cmd_valid),
    .i_icb_cmd_ready        (icb_cmd_ready),
    .i_icb_cmd_read         (icb_cmd_read ),
    .i_icb_cmd_addr         (icb_cmd_addr ),
    .i_icb_cmd_wdata        (icb_cmd_wdata),
    .i_icb_cmd_wmask        (icb_cmd_wmask),
    .i_icb_cmd_lock         (icb_cmd_lock),
    .i_icb_cmd_excl         (icb_cmd_excl),
    .i_icb_cmd_size         (icb_cmd_size ),
    .i_icb_cmd_beat         (icb_cmd_beat),
    .i_icb_cmd_xlen         (icb_cmd_xlen  ),
    .i_icb_cmd_xburst       (icb_cmd_xburst),
    .i_icb_cmd_modes        (icb_cmd_modes ),
    .i_icb_cmd_dmode        (icb_cmd_dmode ),
    .i_icb_cmd_attri        (icb_cmd_attri ),
    .i_icb_rsp_valid        (icb_rsp_valid),
    .i_icb_rsp_ready        (icb_rsp_ready),
    .i_icb_rsp_err          (icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (icb_rsp_rdata),
    .i_icb_cmd_usr          (icb_cmd_usr),
    .i_icb_rsp_usr          (icb_rsp_usr),
    .o_icb_cmd_usr          (buf_icb_cmd_usr),
    .o_icb_rsp_usr          (buf_icb_rsp_usr),
    .o_icb_cmd_sel          (),
    .o_icb_cmd_valid        (buf_icb_cmd_valid),
    .o_icb_cmd_ready        (buf_icb_cmd_ready),
    .o_icb_cmd_read         (buf_icb_cmd_read ),
    .o_icb_cmd_addr         (buf_icb_cmd_addr ),
    .o_icb_cmd_wdata        (buf_icb_cmd_wdata),
    .o_icb_cmd_wmask        (buf_icb_cmd_wmask),
    .o_icb_cmd_lock         (buf_icb_cmd_lock ),
    .o_icb_cmd_size         (buf_icb_cmd_size ),
    .o_icb_cmd_beat         (buf_icb_cmd_beat  ),
    .o_icb_cmd_excl         (buf_icb_cmd_excl  ),
    .o_icb_cmd_xlen         (buf_icb_cmd_xlen  ),
    .o_icb_cmd_xburst       (buf_icb_cmd_xburst),
    .o_icb_cmd_modes        (buf_icb_cmd_modes ),
    .o_icb_cmd_dmode        (buf_icb_cmd_dmode ),
    .o_icb_cmd_attri        (buf_icb_cmd_attri ),
    .o_icb_rsp_valid        (buf_icb_rsp_valid),
    .o_icb_rsp_ready        (buf_icb_rsp_ready),
    .o_icb_rsp_err          (buf_icb_rsp_err  ),
    .o_icb_rsp_rdata        (buf_icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (buf_icb_rsp_excl_ok),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
  wire pend_active;
  e603_subsys_gnrl_usr_ficb2ahbl
  #(
    .CMD_UW(CMD_UW),
    .RSP_UW(RSP_UW),
      .MON_DATA_WIDTH(MON_DATA_WIDTH),
      .AW(AW),
      .DW(DW)
    ) u_icb2ahbl(
    .bus_clk_en        (ratio_ahbl_clk_en),
    .icb2ahbl_pend_active(pend_active),
    .icb_cmd_sel       (buf_icb_cmd_valid   ),
    .icb_cmd_valid     (buf_icb_cmd_valid),
    .icb_cmd_ready     (buf_icb_cmd_ready),
    .icb_cmd_read      (buf_icb_cmd_read ),
    .icb_cmd_addr      (buf_icb_cmd_addr ),
    .icb_cmd_wdata     (buf_icb_cmd_wdata),
    .icb_cmd_wmask     (buf_icb_cmd_wmask),
    .icb_cmd_size      (buf_icb_cmd_size ),
    .icb_cmd_lock      (buf_icb_cmd_lock ),
    .icb_cmd_excl      (buf_icb_cmd_excl),
    .icb_cmd_beat      (buf_icb_cmd_beat  ),
    .icb_cmd_xlen      (buf_icb_cmd_xlen  ),
    .icb_cmd_xburst    (buf_icb_cmd_xburst),
    .icb_cmd_modes     (buf_icb_cmd_modes ),
    .icb_cmd_dmode     (buf_icb_cmd_dmode ),
    .icb_cmd_attri     (buf_icb_cmd_attri ),
    .icb_rsp_valid     (buf_icb_rsp_valid),
    .icb_rsp_ready     (buf_icb_rsp_ready),
    .icb_rsp_err       (buf_icb_rsp_err  ),
    .icb_rsp_rdata     (buf_icb_rsp_rdata),
    .icb_rsp_excl_ok   (buf_icb_rsp_excl_ok),
    .ahbl_htrans       (ratio_htrans  ),
    .ahbl_hwrite       (ratio_hwrite  ),
    .ahbl_haddr        (ratio_haddr   ),
    .ahbl_hsize        (ratio_hsize   ),
    .ahbl_hmastlock    (ratio_hmastlock   ),
    .ahbl_hburst       (ratio_hburst  ),
    .ahbl_hwdata       (ratio_hwdata  ),
    .ahbl_hprot        (ratio_hprot   ),
    .ahbl_hrdata       (ratio_hrdata  ),
    .ahbl_hresp        (ratio_hresp   ),
    .ahbl_hready       (ratio_hready  ),
    .ahbl_hexcl        (),
    .ahbl_hattri       (),
    .ahbl_master       (),
    .ahbl_hresp_exok   (1'b0),
    .ahbl_huser        (ratio_huser   ),
    .icb_cmd_usr      (buf_icb_cmd_usr ),
    .icb_rsp_usr      (buf_icb_rsp_usr ),
    .ahbl_hruser       (ratio_hruser   ),
    .clk               (clk  ),
    .rst_n             (rst_n)
  );
  assign icb2ahbl_ratio_active = pend_active | buffer_active;
  assign icb2ahbl_pend_active = pend_active;
endmodule
module e603_subsys_gnrl_usr_ficb2ahbl_async # (
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter OUTS_CNT_W = 4,
  parameter MON_DATA_WIDTH = 2,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 1,
  parameter ASYNC_FIFO_DP = 4,
  parameter ASYNC_FIFO_DP_PTR_W = 2,
  parameter AW = 32,
  parameter DW = 32
)(
  output icb2ahbl_async_icb_active,
  output icb2ahbl_async_ahbl_active,
  output icb2ahbl_pend_active,
  input  icb_clk,
  input  icb_rst_n,
  input  async_ahbl_clk,
  input  async_ahbl_rst_n,
  input  [CMD_UW -1:0] icb_cmd_usr,
  output [RSP_UW -1:0] icb_rsp_usr,
  output [CMD_UW              -1:0] async_huser,
  input  [RSP_UW              -1:0] async_hruser,
  input             icb_cmd_valid,
  output            icb_cmd_ready,
  input  [AW-1:0]   icb_cmd_addr,
  input             icb_cmd_read,
  input  [DW-1:0]   icb_cmd_wdata,
  input  [DW/8-1:0] icb_cmd_wmask,
  input  [2:0]      icb_cmd_size,
  input             icb_cmd_sel,
  input             icb_cmd_lock,
  input             icb_cmd_excl,
  input  [1:0]      icb_cmd_beat,
  input  [7:0]      icb_cmd_xlen,
  input  [1:0]      icb_cmd_xburst,
  input  [1:0]      icb_cmd_modes,
  input             icb_cmd_dmode,
  input  [2:0]      icb_cmd_attri,
  output            icb_rsp_valid,
  input             icb_rsp_ready,
  output            icb_rsp_err,
  output            icb_rsp_excl_ok,
  output [DW-1:0]   icb_rsp_rdata,
  output [1:0]      async_htrans,
  output            async_hwrite,
  output            async_hmastlock,
  output [2:0]      async_hsize,
  output [2:0]      async_hburst,
  output [3:0]      async_hprot,
  output [DW-1:0]   async_hwdata,
  output [AW-1:0]   async_haddr,
  input  [DW-1:0]   async_hrdata,
  input  [1:0]      async_hresp,
  input             async_hready
  );
  wire icb2icb_async_i_active;
  wire icb2icb_async_o_active;
  wire            async_icb_cmd_valid;
  wire            async_icb_cmd_ready;
  wire [AW-1:0]   async_icb_cmd_addr;
  wire            async_icb_cmd_read;
  wire [DW-1:0]   async_icb_cmd_wdata;
  wire [DW/8-1:0] async_icb_cmd_wmask;
  wire [2:0]      async_icb_cmd_size;
  wire            async_icb_cmd_sel;
  wire            async_icb_cmd_lock;
  wire            async_icb_cmd_excl;
  wire  [1:0]     async_icb_cmd_beat;
  wire  [7:0]     async_icb_cmd_xlen;
  wire  [1:0]     async_icb_cmd_xburst;
  wire  [1:0]     async_icb_cmd_modes;
  wire            async_icb_cmd_dmode;
  wire  [2:0]     async_icb_cmd_attri;
  wire            async_icb_rsp_valid;
  wire            async_icb_rsp_ready;
  wire            async_icb_rsp_err  ;
  wire            async_icb_rsp_excl_ok  ;
  wire [DW-1:0]   async_icb_rsp_rdata;
  wire [CMD_UW-1:0]   async_icb_cmd_usr;
  wire [RSP_UW-1:0]   async_icb_rsp_usr;
  wire [CMD_UW-1:0]   o_icb_cmd_usr;
  wire [RSP_UW-1:0]   o_icb_rsp_usr;
  wire            o_icb_cmd_valid;
  wire            o_icb_cmd_ready;
  wire [AW-1:0]   o_icb_cmd_addr;
  wire            o_icb_cmd_read;
  wire [DW-1:0]   o_icb_cmd_wdata;
  wire [DW/8-1:0] o_icb_cmd_wmask;
  wire [2:0]      o_icb_cmd_size;
  wire            o_icb_cmd_sel;
  wire            o_icb_cmd_lock;
  wire            o_icb_cmd_excl;
  wire  [1:0]     o_icb_cmd_beat;
  wire  [7:0]     o_icb_cmd_xlen;
  wire  [1:0]     o_icb_cmd_xburst;
  wire  [1:0]     o_icb_cmd_modes;
  wire            o_icb_cmd_dmode;
  wire  [2:0]     o_icb_cmd_attri;
  wire            o_icb_rsp_valid;
  wire            o_icb_rsp_ready;
  wire            o_icb_rsp_err  ;
  wire            o_icb_rsp_excl_ok  ;
  wire [DW-1:0]   o_icb_rsp_rdata;
  e603_subsys_gnrl_ficb_async # (
    .RSP_ALWAYS_READY(0),
    .OUTS_CNT_W(OUTS_CNT_W),
    .SYNC_DP (SYNC_DP),
    .ASYNC_FIFO   (ASYNC_FIFO   ),
    .ASYNC_FIFO_DP(ASYNC_FIFO_DP),
    .ASYNC_FIFO_DP_PTR_W(ASYNC_FIFO_DP_PTR_W),
    .AW    (AW),
    .DW    (DW),
    .CMD_UW (CMD_UW),
    .RSP_UW (RSP_UW)
  )u_icb2icb_async(
    .icb2icb_async_i_active   (icb2icb_async_i_active),
    .icb2icb_async_o_active   (icb2icb_async_o_active),
    .i_clk                  (icb_clk),
    .i_rst_n                (icb_rst_n),
    .i_icb_cmd_sel          (icb_cmd_sel),
    .i_icb_cmd_valid        (icb_cmd_valid),
    .i_icb_cmd_ready        (icb_cmd_ready),
    .i_icb_cmd_read         (icb_cmd_read ),
    .i_icb_cmd_addr         (icb_cmd_addr ),
    .i_icb_cmd_wdata        (icb_cmd_wdata),
    .i_icb_cmd_wmask        (icb_cmd_wmask),
    .i_icb_cmd_lock         (icb_cmd_lock ),
    .i_icb_cmd_excl         (icb_cmd_excl ),
    .i_icb_cmd_size         (icb_cmd_size ),
    .i_icb_cmd_beat         (icb_cmd_beat),
    .i_icb_cmd_xlen         (icb_cmd_xlen  ),
    .i_icb_cmd_xburst       (icb_cmd_xburst),
    .i_icb_cmd_modes        (icb_cmd_modes ),
    .i_icb_cmd_dmode        (icb_cmd_dmode ),
    .i_icb_cmd_attri        (icb_cmd_attri ),
    .i_icb_rsp_valid        (icb_rsp_valid),
    .i_icb_rsp_ready        (icb_rsp_ready),
    .i_icb_rsp_err          (icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (icb_rsp_rdata),
    .i_icb_cmd_usr          (icb_cmd_usr),
    .i_icb_rsp_usr          (icb_rsp_usr),
    .o_icb_cmd_usr          (async_icb_cmd_usr),
    .o_icb_rsp_usr          (async_icb_rsp_usr),
    .o_clk                  (async_ahbl_clk),
    .o_rst_n                (async_ahbl_rst_n),
    .o_icb_cmd_sel       (),
    .o_icb_cmd_valid     (async_icb_cmd_valid),
    .o_icb_cmd_ready     (async_icb_cmd_ready),
    .o_icb_cmd_read      (async_icb_cmd_read ),
    .o_icb_cmd_addr      (async_icb_cmd_addr ),
    .o_icb_cmd_wdata     (async_icb_cmd_wdata),
    .o_icb_cmd_wmask     (async_icb_cmd_wmask),
    .o_icb_cmd_size      (async_icb_cmd_size ),
    .o_icb_cmd_beat      (async_icb_cmd_beat  ),
    .o_icb_cmd_lock      (async_icb_cmd_lock  ),
    .o_icb_cmd_excl      (async_icb_cmd_excl  ),
    .o_icb_cmd_xlen      (async_icb_cmd_xlen  ),
    .o_icb_cmd_xburst    (async_icb_cmd_xburst),
    .o_icb_cmd_modes     (async_icb_cmd_modes ),
    .o_icb_cmd_dmode     (async_icb_cmd_dmode ),
    .o_icb_cmd_attri     (async_icb_cmd_attri ),
    .o_icb_rsp_valid        (async_icb_rsp_valid),
    .o_icb_rsp_ready        (async_icb_rsp_ready),
    .o_icb_rsp_err          (async_icb_rsp_err  ),
    .o_icb_rsp_rdata        (async_icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (async_icb_rsp_excl_ok) 
  );
  wire o_buffer_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(0),
    .O_SUPPORT_RATIO(0),
    .AW    (AW),
    .DW    (DW),
    .CMD_DP(0),
    .RSP_BYPBUF(1),
    .RSP_DP(2),
    .OUTS_CNT_W   (2),
    .RSP_ALWAYS_READY(1),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .CMD_UW (CMD_UW),
    .RSP_UW (RSP_UW)
  )u_icb_buffer(
    .i_clk_en (1'b1),
    .o_clk_en (1'b1),
    .icb_buffer_active      (o_buffer_active),
    .i_icb_cmd_sel          (async_icb_cmd_valid),
    .i_icb_cmd_valid        (async_icb_cmd_valid),
    .i_icb_cmd_ready        (async_icb_cmd_ready),
    .i_icb_cmd_read         (async_icb_cmd_read ),
    .i_icb_cmd_addr         (async_icb_cmd_addr ),
    .i_icb_cmd_wdata        (async_icb_cmd_wdata),
    .i_icb_cmd_wmask        (async_icb_cmd_wmask),
    .i_icb_cmd_lock         (async_icb_cmd_lock ),
    .i_icb_cmd_excl         (async_icb_cmd_excl ),
    .i_icb_cmd_size         (async_icb_cmd_size ),
    .i_icb_cmd_beat         (async_icb_cmd_beat),
    .i_icb_cmd_xlen         (async_icb_cmd_xlen  ),
    .i_icb_cmd_xburst       (async_icb_cmd_xburst),
    .i_icb_cmd_modes        (async_icb_cmd_modes ),
    .i_icb_cmd_dmode        (async_icb_cmd_dmode ),
    .i_icb_cmd_attri        (async_icb_cmd_attri ),
    .i_icb_rsp_valid        (async_icb_rsp_valid),
    .i_icb_rsp_ready        (async_icb_rsp_ready),
    .i_icb_rsp_err          (async_icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (async_icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (async_icb_rsp_rdata),
    .i_icb_cmd_usr          (async_icb_cmd_usr),
    .i_icb_rsp_usr          (async_icb_rsp_usr),
    .o_icb_cmd_usr          (o_icb_cmd_usr),
    .o_icb_rsp_usr          (o_icb_rsp_usr),
    .o_icb_cmd_sel          (),
    .o_icb_cmd_valid        (o_icb_cmd_valid),
    .o_icb_cmd_ready        (o_icb_cmd_ready),
    .o_icb_cmd_read         (o_icb_cmd_read ),
    .o_icb_cmd_addr         (o_icb_cmd_addr ),
    .o_icb_cmd_wdata        (o_icb_cmd_wdata),
    .o_icb_cmd_wmask        (o_icb_cmd_wmask),
    .o_icb_cmd_lock         (o_icb_cmd_lock ),
    .o_icb_cmd_size         (o_icb_cmd_size ),
    .o_icb_cmd_beat         (o_icb_cmd_beat  ),
    .o_icb_cmd_excl         (o_icb_cmd_excl  ),
    .o_icb_cmd_xlen         (o_icb_cmd_xlen  ),
    .o_icb_cmd_xburst       (o_icb_cmd_xburst),
    .o_icb_cmd_modes        (o_icb_cmd_modes ),
    .o_icb_cmd_dmode        (o_icb_cmd_dmode ),
    .o_icb_cmd_attri        (o_icb_cmd_attri ),
    .o_icb_rsp_valid        (o_icb_rsp_valid),
    .o_icb_rsp_ready        (o_icb_rsp_ready),
    .o_icb_rsp_err          (o_icb_rsp_err  ),
    .o_icb_rsp_rdata        (o_icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (o_icb_rsp_excl_ok),
    .clk   (async_ahbl_clk  ),
    .rst_n (async_ahbl_rst_n)
  );
  wire icb2ahbl_pend_active_ahbclk;
  e603_subsys_gnrl_usr_ficb2ahbl
  #(
    .CMD_UW(CMD_UW),
    .RSP_UW(RSP_UW),
      .MON_DATA_WIDTH(MON_DATA_WIDTH),
      .AW(AW),
      .DW(DW)
    ) u_icb2ahbl(
    .bus_clk_en        (1'b1),
    .icb2ahbl_pend_active(icb2ahbl_pend_active_ahbclk),
    .icb_cmd_sel       (o_icb_cmd_valid),
    .icb_cmd_valid     (o_icb_cmd_valid),
    .icb_cmd_ready     (o_icb_cmd_ready),
    .icb_cmd_read      (o_icb_cmd_read ),
    .icb_cmd_addr      (o_icb_cmd_addr ),
    .icb_cmd_wdata     (o_icb_cmd_wdata),
    .icb_cmd_wmask     (o_icb_cmd_wmask),
    .icb_cmd_size      (o_icb_cmd_size ),
    .icb_cmd_beat      (o_icb_cmd_beat  ),
    .icb_cmd_lock      (o_icb_cmd_lock  ),
    .icb_cmd_excl      (o_icb_cmd_excl  ),
    .icb_cmd_xlen      (o_icb_cmd_xlen  ),
    .icb_cmd_xburst    (o_icb_cmd_xburst),
    .icb_cmd_modes     (o_icb_cmd_modes ),
    .icb_cmd_dmode     (o_icb_cmd_dmode ),
    .icb_cmd_attri     (o_icb_cmd_attri ),
    .icb_rsp_valid     (o_icb_rsp_valid),
    .icb_rsp_ready     (o_icb_rsp_ready),
    .icb_rsp_err       (o_icb_rsp_err  ),
    .icb_rsp_rdata     (o_icb_rsp_rdata),
    .icb_rsp_excl_ok   (o_icb_rsp_excl_ok),
    .ahbl_htrans       (async_htrans  ),
    .ahbl_hwrite       (async_hwrite  ),
    .ahbl_haddr        (async_haddr   ),
    .ahbl_hsize        (async_hsize   ),
    .ahbl_hmastlock    (async_hmastlock   ),
    .ahbl_hburst       (async_hburst  ),
    .ahbl_hwdata       (async_hwdata  ),
    .ahbl_hprot        (async_hprot   ),
    .ahbl_hrdata       (async_hrdata  ),
    .ahbl_hresp        (async_hresp   ),
    .ahbl_hready       (async_hready  ),
    .ahbl_hexcl        (),
    .ahbl_hattri       (),
    .ahbl_master       (),
    .ahbl_hresp_exok   (1'b0),
    .icb_cmd_usr      (o_icb_cmd_usr ),
    .icb_rsp_usr      (o_icb_rsp_usr ),
    .ahbl_huser        (async_huser   ),
    .ahbl_hruser       (async_hruser   ),
    .clk   (async_ahbl_clk  ),
    .rst_n (async_ahbl_rst_n)
  );
 assign icb2ahbl_async_icb_active = icb2icb_async_i_active;
 assign icb2ahbl_async_ahbl_active = icb2icb_async_o_active | icb2ahbl_pend_active_ahbclk | o_buffer_active;
 assign icb2ahbl_pend_active = 1'b0;
endmodule
module e603_subsys_gnrl_usr_ahbl2ficb_ratio #(
    parameter SUPPORT_ICB_BURST = 0,
    parameter OUTS_CNT_W = 4,
    parameter SUPPORT_RATIO = 0,
    parameter CMD_DP = 0,
    parameter RSP_DP = 0,
    parameter RSP_BYPBUF = 0,
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter WR_EARLY_RETURN = 1,
    parameter AW = 32,
    parameter DW = 32
)(
  output ahbl2icb_ratio_active,
  input  icb_clk_en,
  input  ratio_ahbl_clk_en,
  input  [1:0]                      ahbl_htrans,
  input                             ahbl_hwrite,
  input                             ahbl_hmastlock,
  input  [2:0]                      ahbl_hsize,
  input  [2:0]                      ahbl_hburst,
  input  [3:0]                      ahbl_hprot,
  input  [DW                  -1:0] ahbl_hwdata,
  input  [AW                  -1:0] ahbl_haddr,
  output [DW                  -1:0] ahbl_hrdata,
  output [1:0]                      ahbl_hresp,
  output                            ahbl_hready,
  output                         icb_cmd_valid,
  input                          icb_cmd_ready,
  output [             AW-1:0]   icb_cmd_addr,
  output                         icb_cmd_read,
  output [        DW-1:0]        icb_cmd_wdata,
  output [        DW/8-1:0]      icb_cmd_wmask,
  output                         icb_cmd_lock,
  output                         icb_cmd_excl,
  output [2:0]                   icb_cmd_size,
  output                         icb_cmd_sel,
  output [1:0]                   icb_cmd_beat,
  output [7:0]                   icb_cmd_xlen,
  output [1:0]                   icb_cmd_xburst,
  output [1:0]                   icb_cmd_modes,
  output                         icb_cmd_dmode,
  output [2:0]                   icb_cmd_attri,
  input                          icb_rsp_valid,
  output                         icb_rsp_ready,
  input                          icb_rsp_err  ,
  input                          icb_rsp_excl_ok,
  input  [        DW-1:0]        icb_rsp_rdata,
  input  [CMD_UW              -1:0] ahbl_huser,
  output [RSP_UW              -1:0] ahbl_hruser,
  output [         RSP_UW-1:0]   icb_cmd_usr,
  input  [        RSP_UW-1:0]    icb_rsp_usr,
  input  clk,
  input  rst_n
  );
  wire ahbl2icb_active;
  wire            buf_icb_cmd_valid;
  wire            buf_icb_cmd_ready;
  wire [AW-1:0]   buf_icb_cmd_addr;
  wire            buf_icb_cmd_read;
  wire  [1:0]     buf_icb_cmd_beat;
  wire  [7:0]     buf_icb_cmd_xlen;
  wire  [1:0]     buf_icb_cmd_xburst;
  wire  [1:0]     buf_icb_cmd_modes;
  wire            buf_icb_cmd_dmode;
  wire  [2:0]     buf_icb_cmd_attri;
  wire [CMD_UW-1:0]   buf_icb_cmd_usr;
  wire [RSP_UW-1:0]   buf_icb_rsp_usr;
  wire [DW-1:0]   buf_icb_cmd_wdata;
  wire [DW/8-1:0] buf_icb_cmd_wmask;
  wire            buf_icb_cmd_lock;
  wire            buf_icb_cmd_excl;
  wire [2:0]      buf_icb_cmd_size;
  wire            buf_icb_rsp_valid;
  wire            buf_icb_rsp_ready;
  wire            buf_icb_rsp_err  ;
  wire            buf_icb_rsp_excl_ok  ;
  wire [DW-1:0]   buf_icb_rsp_rdata;
  e603_subsys_gnrl_usr_ahbl2ficb
  #(
      .SUPPORT_ICB_BURST(SUPPORT_ICB_BURST),
      .OUTS_CNT_W(OUTS_CNT_W),
      .CMD_UW(CMD_UW),
      .RSP_UW(RSP_UW),
      .WR_EARLY_RETURN(WR_EARLY_RETURN),
      .AW(AW),
      .DW(DW)
    ) u_ahbl2icb(
    .bus_clk_en        (ratio_ahbl_clk_en),
    .ahbl2icb_active   (ahbl2icb_active),
    .icb_cmd_sel       (),
    .icb_cmd_valid     (buf_icb_cmd_valid),
    .icb_cmd_ready     (buf_icb_cmd_ready),
    .icb_cmd_read      (buf_icb_cmd_read ),
    .icb_cmd_addr      (buf_icb_cmd_addr ),
    .icb_cmd_wdata     (buf_icb_cmd_wdata),
    .icb_cmd_wmask     (buf_icb_cmd_wmask),
    .icb_cmd_size      (buf_icb_cmd_size ),
    .icb_cmd_lock      (buf_icb_cmd_lock ),
    .icb_cmd_excl      (buf_icb_cmd_excl),
    .icb_cmd_beat      (buf_icb_cmd_beat  ),
    .icb_cmd_xlen      (buf_icb_cmd_xlen  ),
    .icb_cmd_xburst    (buf_icb_cmd_xburst),
    .icb_cmd_modes     (buf_icb_cmd_modes ),
    .icb_cmd_dmode     (buf_icb_cmd_dmode ),
    .icb_cmd_attri     (buf_icb_cmd_attri ),
    .icb_cmd_usr       (buf_icb_cmd_usr),
    .icb_rsp_usr       (buf_icb_rsp_usr),
        .ahbl_huser      (ahbl_huser),
        .ahbl_hruser      (ahbl_hruser),
    .icb_rsp_valid     (buf_icb_rsp_valid),
    .icb_rsp_ready     (buf_icb_rsp_ready),
    .icb_rsp_err       (buf_icb_rsp_err  ),
    .icb_rsp_rdata     (buf_icb_rsp_rdata),
    .icb_rsp_excl_ok   (buf_icb_rsp_excl_ok),
    .ahbl_hsel       (1'b1      ),
    .ahbl_htrans     (ahbl_htrans    ),
    .ahbl_hwrite     (ahbl_hwrite    ),
    .ahbl_haddr      (ahbl_haddr     ),
    .ahbl_hsize      (ahbl_hsize     ),
    .ahbl_hprot      (ahbl_hprot      ),
    .ahbl_hwdata     (ahbl_hwdata    ),
    .ahbl_hmastlock  (ahbl_hmastlock ),
    .ahbl_hburst     (ahbl_hburst),
    .ahbl_hexcl      (1'b0),
    .ahbl_hrdata     (ahbl_hrdata    ),
    .ahbl_hresp      (ahbl_hresp     ),
    .ahbl_hready_in  (ahbl_hready),
    .ahbl_hready_out (ahbl_hready),
    .ahbl_hresp_exok (),
    .clk               (clk  ),
    .rst_n             (rst_n)
  );
  wire buffer_active;
  e603_subsys_gnrl_ficb_buffer # (
    .I_SUPPORT_RATIO(SUPPORT_RATIO),
    .O_SUPPORT_RATIO(SUPPORT_RATIO),
    .OUTS_CNT_W   (OUTS_CNT_W),
    .AW    (AW),
    .DW    (DW),
    .CMD_DP(CMD_DP),
    .RSP_DP(RSP_DP),
    .RSP_BYPBUF(RSP_BYPBUF),
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .RSP_ALWAYS_READY(0),
    .CMD_UW (CMD_UW
            ),
    .RSP_UW (RSP_UW)
  )u_icb_buffer(
    .i_clk_en (ratio_ahbl_clk_en),
    .o_clk_en (icb_clk_en),
    .icb_buffer_active      (buffer_active),
    .i_icb_cmd_sel          (buf_icb_cmd_valid),
    .i_icb_cmd_valid        (buf_icb_cmd_valid),
    .i_icb_cmd_ready        (buf_icb_cmd_ready),
    .i_icb_cmd_read         (buf_icb_cmd_read ),
    .i_icb_cmd_addr         (buf_icb_cmd_addr ),
    .i_icb_cmd_wdata        (buf_icb_cmd_wdata),
    .i_icb_cmd_wmask        (buf_icb_cmd_wmask),
    .i_icb_cmd_lock         (buf_icb_cmd_lock ),
    .i_icb_cmd_excl         (buf_icb_cmd_excl ),
    .i_icb_cmd_size         (buf_icb_cmd_size ),
    .i_icb_cmd_beat         (buf_icb_cmd_beat  ),
    .i_icb_cmd_xlen         (buf_icb_cmd_xlen  ),
    .i_icb_cmd_xburst       (buf_icb_cmd_xburst),
    .i_icb_cmd_modes        (buf_icb_cmd_modes ),
    .i_icb_cmd_dmode        (buf_icb_cmd_dmode ),
    .i_icb_cmd_attri        (buf_icb_cmd_attri ),
    .i_icb_cmd_usr          ({buf_icb_cmd_usr
                             }),
    .i_icb_rsp_usr          (buf_icb_rsp_usr),
    .o_icb_cmd_usr          ({icb_cmd_usr
                             }),
    .o_icb_rsp_usr          (icb_rsp_usr  ),
    .i_icb_rsp_valid        (buf_icb_rsp_valid),
    .i_icb_rsp_ready        (buf_icb_rsp_ready),
    .i_icb_rsp_err          (buf_icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (buf_icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (buf_icb_rsp_rdata),
    .o_icb_cmd_sel          (icb_cmd_sel  ),
    .o_icb_cmd_valid        (icb_cmd_valid),
    .o_icb_cmd_ready        (icb_cmd_ready),
    .o_icb_cmd_read         (icb_cmd_read ),
    .o_icb_cmd_addr         (icb_cmd_addr ),
    .o_icb_cmd_wdata        (icb_cmd_wdata),
    .o_icb_cmd_wmask        (icb_cmd_wmask),
    .o_icb_cmd_lock         (icb_cmd_lock ),
    .o_icb_cmd_size         (icb_cmd_size ),
    .o_icb_cmd_beat         (icb_cmd_beat  ),
    .o_icb_cmd_excl         (icb_cmd_excl  ),
    .o_icb_cmd_xlen         (icb_cmd_xlen  ),
    .o_icb_cmd_xburst       (icb_cmd_xburst),
    .o_icb_cmd_modes        (icb_cmd_modes ),
    .o_icb_cmd_dmode        (icb_cmd_dmode ),
    .o_icb_cmd_attri        (icb_cmd_attri ),
    .o_icb_rsp_valid        (icb_rsp_valid),
    .o_icb_rsp_ready        (icb_rsp_ready),
    .o_icb_rsp_err          (icb_rsp_err  ),
    .o_icb_rsp_rdata        (icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (icb_rsp_excl_ok),
    .clk                    (clk  ),
    .rst_n                  (rst_n)
  );
  assign ahbl2icb_ratio_active = ahbl2icb_active | buffer_active;
endmodule
module e603_subsys_gnrl_usr_ahbl2ficb_async # (
    parameter SUPPORT_ICB_BURST = 0,
    parameter OUTS_CNT_W = 4,
    parameter CMD_UW = 1,
    parameter RSP_UW = 1,
    parameter WR_EARLY_RETURN = 1,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 1,
  parameter ASYNC_FIFO_DP = 4,
  parameter ASYNC_FIFO_DP_PTR_W = 2,
  parameter AW = 32,
  parameter DW = 32
)(
  output ahbl2icb_async_ahbl_active,
  output ahbl2icb_async_icb_active,
  input  icb_clk,
  input  icb_rst_n,
  input  async_ahbl_clk,
  input  async_ahbl_rst_n,
  input  [1:0]                      ahbl_htrans,
  input                             ahbl_hwrite,
  input                             ahbl_hmastlock,
  input  [2:0]                      ahbl_hsize,
  input  [2:0]                      ahbl_hburst,
  input  [3:0]                      ahbl_hprot,
  input  [DW                  -1:0] ahbl_hwdata,
  input  [AW                  -1:0] ahbl_haddr,
  output [DW                  -1:0] ahbl_hrdata,
  output [1:0]                      ahbl_hresp,
  output                            ahbl_hready,
  output                         icb_cmd_valid,
  input                          icb_cmd_ready,
  output [             AW-1:0]   icb_cmd_addr,
  output                         icb_cmd_read,
  output [        DW-1:0]        icb_cmd_wdata,
  output [        DW/8-1:0]      icb_cmd_wmask,
  output                         icb_cmd_lock,
  output                         icb_cmd_excl,
  output [2:0]                   icb_cmd_size,
  output                         icb_cmd_sel,
  output [1:0]                   icb_cmd_beat,
  output [7:0]                   icb_cmd_xlen,
  output [1:0]                   icb_cmd_xburst,
  output [1:0]                   icb_cmd_modes,
  output                         icb_cmd_dmode,
  output [2:0]                   icb_cmd_attri,
  input  [CMD_UW              -1:0] ahbl_huser,
  output [RSP_UW              -1:0] ahbl_hruser,
  output [         RSP_UW-1:0]   icb_cmd_usr,
  input  [        RSP_UW-1:0]    icb_rsp_usr,
  input                          icb_rsp_valid,
  output                         icb_rsp_ready,
  input                          icb_rsp_err  ,
  input                          icb_rsp_excl_ok,
  input  [        DW-1:0]        icb_rsp_rdata
  );
  wire icb2icb_async_i_active;
  wire icb2icb_async_o_active;
  wire ahbl2icb_active;
  wire            async_icb_cmd_valid;
  wire            async_icb_cmd_ready;
  wire [AW-1:0]   async_icb_cmd_addr;
  wire            async_icb_cmd_read;
  wire [DW-1:0]   async_icb_cmd_wdata;
  wire [DW/8-1:0] async_icb_cmd_wmask;
  wire [2:0]      async_icb_cmd_size;
  wire            async_icb_cmd_sel;
  wire            async_icb_cmd_lock;
  wire            async_icb_cmd_excl;
  wire  [1:0]     async_icb_cmd_beat;
  wire  [7:0]     async_icb_cmd_xlen;
  wire  [1:0]     async_icb_cmd_xburst;
  wire  [1:0]     async_icb_cmd_modes;
  wire            async_icb_cmd_dmode;
  wire  [2:0]     async_icb_cmd_attri;
  wire            async_icb_rsp_valid;
  wire            async_icb_rsp_ready;
  wire            async_icb_rsp_err  ;
  wire            async_icb_rsp_excl_ok  ;
  wire [DW-1:0]   async_icb_rsp_rdata;
  wire [CMD_UW-1:0]   async_icb_cmd_usr;
  wire [RSP_UW-1:0]   async_icb_rsp_usr;
  e603_subsys_gnrl_usr_ahbl2ficb
  #(
      .SUPPORT_ICB_BURST(SUPPORT_ICB_BURST),
      .OUTS_CNT_W(OUTS_CNT_W),
      .CMD_UW(CMD_UW),
      .RSP_UW(RSP_UW),
      .WR_EARLY_RETURN(WR_EARLY_RETURN),
      .AW(AW),
      .DW(DW)
    ) u_ahbl2icb(
    .bus_clk_en        (1'b1),
    .ahbl2icb_active   (ahbl2icb_active),
    .icb_cmd_sel       (   ),
    .icb_cmd_valid     (async_icb_cmd_valid),
    .icb_cmd_ready     (async_icb_cmd_ready),
    .icb_cmd_read      (async_icb_cmd_read ),
    .icb_cmd_addr      (async_icb_cmd_addr ),
    .icb_cmd_wdata     (async_icb_cmd_wdata),
    .icb_cmd_wmask     (async_icb_cmd_wmask),
    .icb_cmd_size      (async_icb_cmd_size ),
    .icb_cmd_lock      (async_icb_cmd_lock ),
    .icb_cmd_excl      (async_icb_cmd_excl),
    .icb_cmd_beat      (async_icb_cmd_beat  ),
    .icb_cmd_xlen      (async_icb_cmd_xlen  ),
    .icb_cmd_xburst    (async_icb_cmd_xburst),
    .icb_cmd_modes     (async_icb_cmd_modes ),
    .icb_cmd_dmode     (async_icb_cmd_dmode ),
    .icb_cmd_attri     (async_icb_cmd_attri ),
    .icb_rsp_valid     (async_icb_rsp_valid),
    .icb_rsp_ready     (async_icb_rsp_ready),
    .icb_rsp_err       (async_icb_rsp_err  ),
    .icb_rsp_rdata     (async_icb_rsp_rdata),
    .icb_rsp_excl_ok   (async_icb_rsp_excl_ok),
    .icb_cmd_usr       (async_icb_cmd_usr),
    .icb_rsp_usr       (async_icb_rsp_usr),
        .ahbl_huser      (ahbl_huser),
        .ahbl_hruser      (ahbl_hruser),
    .ahbl_hsel       (1'b1      ),
    .ahbl_htrans     (ahbl_htrans    ),
    .ahbl_hwrite     (ahbl_hwrite    ),
    .ahbl_haddr      (ahbl_haddr     ),
    .ahbl_hsize      (ahbl_hsize     ),
    .ahbl_hwdata     (ahbl_hwdata    ),
    .ahbl_hmastlock  (ahbl_hmastlock ),
    .ahbl_hburst     (ahbl_hburst),
    .ahbl_hexcl      (1'b0),
    .ahbl_hprot      (ahbl_hprot      ),
    .ahbl_hrdata     (ahbl_hrdata    ),
    .ahbl_hresp      (ahbl_hresp     ),
    .ahbl_hready_in  (ahbl_hready),
    .ahbl_hready_out (ahbl_hready),
    .ahbl_hresp_exok (),
    .clk               (async_ahbl_clk  ),
    .rst_n             (async_ahbl_rst_n)
  );
  e603_subsys_gnrl_ficb_async # (
    .RSP_ALWAYS_READY(0),
    .OUTS_CNT_W(OUTS_CNT_W),
    .SYNC_DP (SYNC_DP),
    .ASYNC_FIFO (ASYNC_FIFO),
    .ASYNC_FIFO_DP(ASYNC_FIFO_DP),
    .ASYNC_FIFO_DP_PTR_W(ASYNC_FIFO_DP_PTR_W),
    .AW    (AW),
    .DW    (DW),
    .CMD_UW (CMD_UW
            ),
    .RSP_UW (RSP_UW)
  )u_icb2icb_async(
    .icb2icb_async_i_active   (icb2icb_async_i_active),
    .icb2icb_async_o_active   (icb2icb_async_o_active),
    .i_clk                  (async_ahbl_clk),
    .i_rst_n                (async_ahbl_rst_n),
    .o_clk                  (icb_clk),
    .o_rst_n                (icb_rst_n),
    .i_icb_cmd_sel          (async_icb_cmd_valid),
    .i_icb_cmd_valid        (async_icb_cmd_valid),
    .i_icb_cmd_ready        (async_icb_cmd_ready),
    .i_icb_cmd_read         (async_icb_cmd_read ),
    .i_icb_cmd_addr         (async_icb_cmd_addr ),
    .i_icb_cmd_wdata        (async_icb_cmd_wdata),
    .i_icb_cmd_wmask        (async_icb_cmd_wmask),
    .i_icb_cmd_lock         (async_icb_cmd_lock   ),
    .i_icb_cmd_excl         (async_icb_cmd_excl   ),
    .i_icb_cmd_size         (async_icb_cmd_size   ),
    .i_icb_cmd_beat         (async_icb_cmd_beat   ),
    .i_icb_cmd_xlen         (async_icb_cmd_xlen   ),
    .i_icb_cmd_xburst       (async_icb_cmd_xburst ),
    .i_icb_cmd_modes        (async_icb_cmd_modes ),
    .i_icb_cmd_dmode        (async_icb_cmd_dmode ),
    .i_icb_cmd_attri        (async_icb_cmd_attri ),
    .i_icb_rsp_valid        (async_icb_rsp_valid),
    .i_icb_rsp_ready        (async_icb_rsp_ready),
    .i_icb_rsp_err          (async_icb_rsp_err  ),
    .i_icb_rsp_excl_ok      (async_icb_rsp_excl_ok),
    .i_icb_rsp_rdata        (async_icb_rsp_rdata),
    .i_icb_cmd_usr          ({async_icb_cmd_usr
                             }),
    .i_icb_rsp_usr          (async_icb_rsp_usr),
    .o_icb_cmd_usr          ({icb_cmd_usr
                             }),
    .o_icb_rsp_usr          (icb_rsp_usr  ),
    .o_icb_cmd_sel       (icb_cmd_sel  ),
    .o_icb_cmd_valid     (icb_cmd_valid),
    .o_icb_cmd_ready     (icb_cmd_ready),
    .o_icb_cmd_read      (icb_cmd_read ),
    .o_icb_cmd_addr      (icb_cmd_addr ),
    .o_icb_cmd_wdata     (icb_cmd_wdata),
    .o_icb_cmd_wmask     (icb_cmd_wmask),
    .o_icb_cmd_size      (icb_cmd_size ),
    .o_icb_cmd_beat      (icb_cmd_beat  ),
    .o_icb_cmd_lock      (icb_cmd_lock  ),
    .o_icb_cmd_excl      (icb_cmd_excl  ),
    .o_icb_cmd_xlen      (icb_cmd_xlen  ),
    .o_icb_cmd_xburst    (icb_cmd_xburst),
    .o_icb_cmd_modes     (icb_cmd_modes ),
    .o_icb_cmd_dmode     (icb_cmd_dmode ),
    .o_icb_cmd_attri     (icb_cmd_attri ),
    .o_icb_rsp_valid        (icb_rsp_valid),
    .o_icb_rsp_ready        (icb_rsp_ready),
    .o_icb_rsp_err          (icb_rsp_err  ),
    .o_icb_rsp_rdata        (icb_rsp_rdata),
    .o_icb_rsp_excl_ok      (icb_rsp_excl_ok) 
  );
 assign ahbl2icb_async_ahbl_active = icb2icb_async_i_active | ahbl2icb_active;
 assign ahbl2icb_async_icb_active = icb2icb_async_o_active;
endmodule
module e603_subsys_gnrl_ficb_rw_splt # (
  parameter ALLOW_DIFF = 1,
  parameter AW = 32,
  parameter DW = 32,
  parameter OUTS_FIFO_DP =4,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr,
  input                         icb_cmd_read,
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]              icb_cmd_wmask,
  input [CMD_UW-1:0]            icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [2:0]                   icb_cmd_size,
  input [7:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]           icb_rsp_usr,
  input                         r_icb_cmd_ready,
  output                        r_icb_cmd_sel,
  output                        r_icb_cmd_valid,
  output[AW-1:0]                r_icb_cmd_addr,
  output                        r_icb_cmd_read,
  output[DW-1:0]                r_icb_cmd_wdata,
  output[DW/8-1:0]              r_icb_cmd_wmask,
  output[CMD_UW-1:0]            r_icb_cmd_usr,
  output[1:0]                   r_icb_cmd_beat,
  output                        r_icb_cmd_lock,
  output                        r_icb_cmd_excl,
  output[2:0]                   r_icb_cmd_size,
  output[7:0]                   r_icb_cmd_xlen,
  output[1:0]                   r_icb_cmd_xburst,
  output[1:0]                   r_icb_cmd_modes,
  output                        r_icb_cmd_dmode,
  output[2:0]                   r_icb_cmd_attri,
  output                        r_icb_rsp_ready,
  input                         r_icb_rsp_valid,
  input                         r_icb_rsp_err  ,
  input                         r_icb_rsp_excl_ok,
  input  [DW-1:0]               r_icb_rsp_rdata,
  input  [RSP_UW-1:0]           r_icb_rsp_usr,
  input                         w_icb_cmd_ready,
  output                        w_icb_cmd_sel,
  output                        w_icb_cmd_valid,
  output[AW-1:0]                w_icb_cmd_addr,
  output                        w_icb_cmd_read,
  output[DW-1:0]                w_icb_cmd_wdata,
  output[DW/8-1:0]              w_icb_cmd_wmask,
  output[CMD_UW-1:0]            w_icb_cmd_usr,
  output[1:0]                   w_icb_cmd_beat,
  output                        w_icb_cmd_lock,
  output                        w_icb_cmd_excl,
  output[2:0]                   w_icb_cmd_size,
  output[7:0]                   w_icb_cmd_xlen,
  output[1:0]                   w_icb_cmd_xburst,
  output[1:0]                   w_icb_cmd_modes,
  output                        w_icb_cmd_dmode,
  output[2:0]                   w_icb_cmd_attri,
  output                        w_icb_rsp_ready,
  input                         w_icb_rsp_valid,
  input                         w_icb_rsp_err  ,
  input                         w_icb_rsp_excl_ok,
  input  [DW-1:0]               w_icb_rsp_rdata,
  input  [RSP_UW-1:0]           w_icb_rsp_usr,
  input                         clk,
  input                         rst_n
  );
   wire [1:0] icb_cmd_splt_indic ={
      (~icb_cmd_read),
      icb_cmd_read
      };
  localparam SPLT_I_NUM = 2;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_sel;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_ready;
  wire [SPLT_I_NUM*AW-1:0] splt_bus_icb_cmd_addr;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_read;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_cmd_wdata;
  wire [SPLT_I_NUM*DW/8-1:0] splt_bus_icb_cmd_wmask;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_beat;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_lock;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_excl;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_size;
  wire [SPLT_I_NUM*CMD_UW-1:0] splt_bus_icb_cmd_usr;
  wire [SPLT_I_NUM*8-1:0] splt_bus_icb_cmd_xlen  ;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_xburst;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_modes ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_dmode ;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_attri ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_ready;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_err;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_excl_ok;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_rsp_rdata;
  wire [SPLT_I_NUM*RSP_UW-1:0] splt_bus_icb_rsp_usr;
  assign {
                             w_icb_cmd_valid,
                             r_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
  assign {
                             w_icb_cmd_sel,
                             r_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
  assign {
                             w_icb_cmd_addr,
                             r_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
  assign {
                             w_icb_cmd_read,
                             r_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
  assign {
                             w_icb_cmd_wdata,
                             r_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
  assign {
                             w_icb_cmd_wmask,
                             r_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
  assign {
                             w_icb_cmd_xburst,
                             r_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
  assign {
                             w_icb_cmd_xlen,
                             r_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
  assign {
                             w_icb_cmd_modes,
                             r_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
  assign {
                             w_icb_cmd_dmode,
                             r_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
  assign {
                             w_icb_cmd_attri,
                             r_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
  assign {
                             w_icb_cmd_beat,
                             r_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
  assign {
                             w_icb_cmd_lock,
                             r_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
  assign {
                             w_icb_cmd_excl,
                             r_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
  assign {
                             w_icb_cmd_size,
                             r_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
  assign {
                             w_icb_cmd_usr,
                             r_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
  assign splt_bus_icb_cmd_ready = {
                             w_icb_cmd_ready,
                             r_icb_cmd_ready
                           };
  assign splt_bus_icb_rsp_valid = {
                             w_icb_rsp_valid,
                             r_icb_rsp_valid
                           };
  assign splt_bus_icb_rsp_err = {
                             w_icb_rsp_err,
                             r_icb_rsp_err
                           };
  assign splt_bus_icb_rsp_excl_ok = {
                             w_icb_rsp_excl_ok,
                             r_icb_rsp_excl_ok
                           };
  assign splt_bus_icb_rsp_rdata = {
                             w_icb_rsp_rdata,
                             r_icb_rsp_rdata
                           };
  assign splt_bus_icb_rsp_usr = {
                             w_icb_rsp_usr,
                             r_icb_rsp_usr
                           };
  assign {
                             w_icb_rsp_ready,
                             r_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
  e603_subsys_gnrl_ficb_splt # (
  .USE_ALL_READY(0),
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (0),
  .FIFO_OUTS_NUM   (OUTS_FIFO_DP),
  .FIFO_CUT_READY  (1),
  .SPLT_NUM   (2),
  .SPLT_PTR_W (2),
  .SPLT_PTR_1HOT (1),
  .CMD_UW     (CMD_UW),
  .RSP_UW     (RSP_UW),
  .AW         (AW),
  .DW         (DW)
  ) u_icb_rw_splt(
  .clk_en(1'b1),
  .splt_active            (),
  .i_icb_splt_indic       (icb_cmd_splt_indic),
  .i_icb_cmd_sel          (icb_cmd_sel )     ,
  .i_icb_cmd_valid        (icb_cmd_valid )     ,
  .i_icb_cmd_ready        (icb_cmd_ready )     ,
  .i_icb_cmd_read         (icb_cmd_read )      ,
  .i_icb_cmd_addr         (icb_cmd_addr )      ,
  .i_icb_cmd_wdata        (icb_cmd_wdata )     ,
  .i_icb_cmd_wmask        (icb_cmd_wmask)      ,
  .i_icb_cmd_beat         (icb_cmd_beat )     ,
  .i_icb_cmd_excl         (icb_cmd_excl )     ,
  .i_icb_cmd_lock         (icb_cmd_lock )     ,
  .i_icb_cmd_size         (icb_cmd_size )     ,
  .i_icb_cmd_xburst       (icb_cmd_xburst),
  .i_icb_cmd_xlen         (icb_cmd_xlen  ),
  .i_icb_cmd_modes        (icb_cmd_modes ),
  .i_icb_cmd_dmode        (icb_cmd_dmode ),
  .i_icb_cmd_attri        (icb_cmd_attri ),
  .i_icb_cmd_usr          (icb_cmd_usr   ),
  .i_icb_rsp_valid        (icb_rsp_valid )     ,
  .i_icb_rsp_ready        (icb_rsp_ready )     ,
  .i_icb_rsp_err          (icb_rsp_err)        ,
  .i_icb_rsp_excl_ok      (icb_rsp_excl_ok)    ,
  .i_icb_rsp_rdata        (icb_rsp_rdata )     ,
  .i_icb_rsp_usr          (icb_rsp_usr )     ,
  .o_bus_icb_cmd_ready    (splt_bus_icb_cmd_ready ) ,
  .o_bus_icb_cmd_valid    (splt_bus_icb_cmd_valid ) ,
  .o_bus_icb_cmd_sel      (splt_bus_icb_cmd_sel   ) ,
  .o_bus_icb_cmd_read     (splt_bus_icb_cmd_read )  ,
  .o_bus_icb_cmd_addr     (splt_bus_icb_cmd_addr )  ,
  .o_bus_icb_cmd_wdata    (splt_bus_icb_cmd_wdata ) ,
  .o_bus_icb_cmd_wmask    (splt_bus_icb_cmd_wmask)  ,
  .o_bus_icb_cmd_beat     (splt_bus_icb_cmd_beat ),
  .o_bus_icb_cmd_excl     (splt_bus_icb_cmd_excl ),
  .o_bus_icb_cmd_lock     (splt_bus_icb_cmd_lock ),
  .o_bus_icb_cmd_size     (splt_bus_icb_cmd_size ),
  .o_bus_icb_cmd_usr      (splt_bus_icb_cmd_usr  ),
  .o_bus_icb_cmd_xburst   (splt_bus_icb_cmd_xburst),
  .o_bus_icb_cmd_xlen     (splt_bus_icb_cmd_xlen  ),
  .o_bus_icb_cmd_modes    (splt_bus_icb_cmd_modes ),
  .o_bus_icb_cmd_dmode    (splt_bus_icb_cmd_dmode ),
  .o_bus_icb_cmd_attri    (splt_bus_icb_cmd_attri ),
  .o_bus_icb_rsp_valid    (splt_bus_icb_rsp_valid ) ,
  .o_bus_icb_rsp_ready    (splt_bus_icb_rsp_ready ) ,
  .o_bus_icb_rsp_err      (splt_bus_icb_rsp_err)    ,
  .o_bus_icb_rsp_excl_ok  (splt_bus_icb_rsp_excl_ok),
  .o_bus_icb_rsp_rdata    (splt_bus_icb_rsp_rdata ) ,
  .o_bus_icb_rsp_usr      (splt_bus_icb_rsp_usr ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
`include "global.v"
module e603_subsys_gnrl_ficb_arbt_id # (
    parameter I_REAL_ID_W = 0,
    parameter ID_W = 4,
  parameter SUPPORT_LOCK = 1,
  parameter PAYLOAD_NORST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter ARBT_SCHEME = 3,
  parameter RRBIN_CUT_TIMING = 0,
  parameter FIFO_OUTS_NUM = 1,
  parameter FIFO_REG_OUT = 0,
  parameter FIFO_CUT_READY = 0,
  parameter ARBT_NUM = 4,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter ARBT_PTR_W = 2
) (
  output             arbt_active,
  input              clk_en,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [DW-1:0]    o_icb_cmd_wdata,
  output [DW/8-1:0]    o_icb_cmd_wmask,
  output [2-1:0]     o_icb_cmd_beat,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [CMD_SIZE_W-1:0]       o_icb_cmd_size,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  output [ID_W-1:0]  o_icb_cmd_id,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0]  o_icb_rsp_id,
  input              o_icb_rsp_last,
  output [ARBT_NUM*1-1:0]     i_bus_icb_cmd_ready,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_valid,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_read,
  input  [ARBT_NUM*AW-1:0]    i_bus_icb_cmd_addr,
  input  [ARBT_NUM*DW-1:0]    i_bus_icb_cmd_wdata,
  input  [ARBT_NUM*DW/8-1:0]    i_bus_icb_cmd_wmask,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_beat ,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_lock ,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_excl ,
  input  [ARBT_NUM*CMD_SIZE_W-1:0]     i_bus_icb_cmd_size ,
  input  [ARBT_NUM*CMD_UW-1:0] i_bus_icb_cmd_usr  ,
  input  [ARBT_NUM*ID_W-1:0]   i_bus_icb_cmd_id  ,
  input  [ARBT_NUM*8-1:0]     i_bus_icb_cmd_xlen,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_xburst,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_modes,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_dmode,
  input  [ARBT_NUM*3-1:0]     i_bus_icb_cmd_attri,
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_valid,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_rsp_ready,
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_err,
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_excl_ok,
  output [ARBT_NUM*DW-1:0]    i_bus_icb_rsp_rdata,
  output [ARBT_NUM*RSP_UW-1:0] i_bus_icb_rsp_usr,
  output [ARBT_NUM*ID_W-1:0] i_bus_icb_rsp_id,
  output [ARBT_NUM     -1:0] i_bus_icb_rsp_last,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_sel_vec,
  input  clk,
  input  rst_n
  );
    localparam I_ICB_IDW_ZERO = (ARBT_NUM > 1) ? ((ID_W == ARBT_PTR_W) ? 1 : 0) : 0;
  localparam ARBT_SCHEME_PRIORITY  = 0;
  localparam ARBT_SCHEME_RROBIN    = 1;
  localparam ARBT_SCHEME_DIRECT_SEL_1HOT = 2;
  localparam ARBT_SCHEME_DIRECT_SEL_PRIORITY = 3;
  localparam ARBT_SCHEME_RROBIN4   = 4;
  localparam ARBT_SCHEME_RROBIN_TIME = 5;
  wire             icb_rsp_valid;
  wire             icb_rsp_ready;
  wire             icb_rsp_err;
  wire             icb_rsp_excl_ok;
  wire [DW-1:0]    icb_rsp_rdata;
  wire [RSP_UW-1:0] icb_rsp_usr;
  wire [ID_W-1:0] icb_rsp_id;
  wire            icb_rsp_last;
  wire [ARBT_PTR_W-1:0] t_icb_rsp_id;
  wire                  t_icb_rsp_last;
  localparam RSP_PACK_W = (2+DW+RSP_UW+ID_W+1);
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata,
                                 o_icb_rsp_id,
                                 o_icb_rsp_last,
                                 o_icb_rsp_usr};
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 icb_rsp_err,
                                 icb_rsp_excl_ok,
                                 icb_rsp_rdata,
                                 icb_rsp_id,
                                 icb_rsp_last,
                                 icb_rsp_usr} = rsp_fifo_o_dat;
      assign rsp_fifo_o_dat = rsp_fifo_i_dat;
      assign icb_rsp_valid = o_icb_rsp_valid;
      assign o_icb_rsp_ready = icb_rsp_ready;
  wire rspid_fifo_empty;
  wire rrobin_active;
  wire rrobin_notime_active;
  wire rrobin_time_active;
  wire rbin4_active;
  wire [ARBT_NUM-1:0] lock_mask_r  ;
  wire [ARBT_NUM-1:0] omask_r;
  wire [ARBT_NUM-1:0] burst_mask_r;
genvar i;
generate 
  if(ARBT_NUM == 1) begin:gen_arbt_num_eq_1
    assign i_bus_icb_cmd_ready = o_icb_cmd_ready    ;
    assign o_icb_cmd_valid     = i_bus_icb_cmd_valid;
    assign o_icb_cmd_sel       = i_bus_icb_cmd_sel_vec  ;
    assign o_icb_cmd_read      = i_bus_icb_cmd_read ;
    assign o_icb_cmd_addr      = i_bus_icb_cmd_addr ;
    assign o_icb_cmd_wdata     = i_bus_icb_cmd_wdata;
    assign o_icb_cmd_wmask     = i_bus_icb_cmd_wmask;
    assign o_icb_cmd_beat      = i_bus_icb_cmd_beat ;
    assign o_icb_cmd_lock      = i_bus_icb_cmd_lock ;
    assign o_icb_cmd_excl      = i_bus_icb_cmd_excl ;
    assign o_icb_cmd_size      = i_bus_icb_cmd_size ;
    assign o_icb_cmd_usr       = i_bus_icb_cmd_usr  ;
    assign o_icb_cmd_id        = i_bus_icb_cmd_id  ;
    assign o_icb_cmd_xlen      = i_bus_icb_cmd_xlen  ;
    assign o_icb_cmd_xburst    = i_bus_icb_cmd_xburst;
    assign o_icb_cmd_modes     = i_bus_icb_cmd_modes ;
    assign o_icb_cmd_dmode     = i_bus_icb_cmd_dmode ;
    assign o_icb_cmd_attri     = i_bus_icb_cmd_attri ;
    assign icb_rsp_ready     = i_bus_icb_rsp_ready;
    assign i_bus_icb_rsp_valid = icb_rsp_valid    ;
    assign i_bus_icb_rsp_err   = icb_rsp_err      ;
    assign i_bus_icb_rsp_excl_ok   = icb_rsp_excl_ok      ;
    assign i_bus_icb_rsp_rdata = icb_rsp_rdata    ;
    assign i_bus_icb_rsp_usr   = icb_rsp_usr      ;
    assign i_bus_icb_rsp_id   = icb_rsp_id      ;
    assign i_bus_icb_rsp_last   = icb_rsp_last      ;
    assign rspid_fifo_empty    = 1'b1;
    assign lock_mask_r = {ARBT_NUM{1'b0}};
    assign omask_r = {ARBT_NUM{1'b0}};
    assign burst_mask_r = {ARBT_NUM{1'b0}};
    assign rbin4_active = 1'b0;
    assign rrobin_active = 1'b0;
    assign rrobin_time_active = 1'b0;
    assign rrobin_notime_active = 1'b0;
  end
  else begin:gen_arbt_num_gt_1
    integer j;
    wire [ARBT_NUM-1:0] i_bus_icb_cmd_grt_vec;
    wire [ARBT_NUM-1:0] i_bus_icb_cmd_sel;
    wire o_icb_cmd_valid_real;
    wire o_icb_cmd_ready_real;
    wire            i_icb_cmd_read [ARBT_NUM-1:0];
    wire [AW-1:0]   i_icb_cmd_addr [ARBT_NUM-1:0];
    wire [DW-1:0]   i_icb_cmd_wdata[ARBT_NUM-1:0];
    wire [DW/8-1:0]   i_icb_cmd_wmask[ARBT_NUM-1:0];
    wire [2-1:0]    i_icb_cmd_beat [ARBT_NUM-1:0];
    wire            i_icb_cmd_lock [ARBT_NUM-1:0];
    wire            i_icb_cmd_excl [ARBT_NUM-1:0];
    wire [CMD_SIZE_W-1:0]    i_icb_cmd_size [ARBT_NUM-1:0];
    wire [CMD_UW-1:0]i_icb_cmd_usr  [ARBT_NUM-1:0];
    wire [ID_W-1:0]i_icb_cmd_id  [ARBT_NUM-1:0];
    wire [7:0]      i_icb_cmd_xlen   [ARBT_NUM-1:0];
    wire [1:0]      i_icb_cmd_xburst [ARBT_NUM-1:0];
    wire [1:0]      i_icb_cmd_modes  [ARBT_NUM-1:0];
    wire            i_icb_cmd_dmode  [ARBT_NUM-1:0];
    wire [2:0]      i_icb_cmd_attri  [ARBT_NUM-1:0];
    reg            sel_o_icb_cmd_read;
    reg [AW-1:0]   sel_o_icb_cmd_addr;
    reg [DW-1:0]   sel_o_icb_cmd_wdata;
    reg [DW/8-1:0]   sel_o_icb_cmd_wmask;
    reg [2-1:0]    sel_o_icb_cmd_beat ;
    reg            sel_o_icb_cmd_lock ;
    reg            sel_o_icb_cmd_excl ;
    reg [CMD_SIZE_W-1:0]    sel_o_icb_cmd_size ;
    reg [CMD_UW-1:0]sel_o_icb_cmd_usr  ;
    reg [ID_W-1:0]sel_o_icb_cmd_id  ;
    reg [7:0]      sel_o_icb_cmd_xlen  ;
    reg [1:0]      sel_o_icb_cmd_xburst;
    reg [1:0]      sel_o_icb_cmd_modes ;
    reg            sel_o_icb_cmd_dmode ;
    reg [2:0]      sel_o_icb_cmd_attri ;
    wire icb_rsp_ready_pre;
    wire icb_rsp_valid_pre;
    wire rspid_fifo_bypass;
    wire rspid_fifo_wen;
    wire rspid_fifo_ren;
    wire rspid_fifo_i_valid;
    wire rspid_fifo_o_valid;
    wire rspid_fifo_i_ready;
    wire rspid_fifo_o_ready;
    wire [ARBT_PTR_W-1:0] rspid_fifo_rdat;
    wire [ARBT_PTR_W-1:0] rspid_fifo_wdat;
    wire rspid_fifo_full;
    reg [ARBT_PTR_W-1:0] i_arbt_indic_id;
    wire [ARBT_NUM*1-1:0] i_bus_icb_cmd_ready_pos;
    wire [ARBT_NUM*1-1:0] i_bus_icb_cmd_valid_pos;
    wire [ARBT_NUM*1-1:0] i_bus_icb_cmd_sel_vec_pos;
    wire arbt_ena;
    wire [ARBT_PTR_W-1:0] icb_rsp_port_id;
    if((ARBT_SCHEME == ARBT_SCHEME_RROBIN) || (ARBT_SCHEME == ARBT_SCHEME_RROBIN_TIME) || (ARBT_SCHEME == ARBT_SCHEME_RROBIN4)) begin: gen_rrobin
        assign omask_r = {ARBT_NUM{1'b0}};
    end
    else begin: gen_not_rrobin
        wire [ARBT_NUM-1:0] omask_nxt;
        wire omask_ena;
        wire omask_set;
        wire omask_clr;
        assign omask_set = o_icb_cmd_valid_real & (~arbt_ena); 
        assign omask_clr = (|omask_r) & (arbt_ena | (~o_icb_cmd_valid_real));
        assign omask_ena = clk_en & (omask_set | omask_clr);
        assign omask_nxt = omask_clr ? {ARBT_NUM{1'b0}} : (~i_bus_icb_cmd_sel); 
e603_subsys_gnrl_dfflr #(ARBT_NUM) omask_dfflr (omask_ena, omask_nxt, omask_r, clk, rst_n);// VPP_NO_REG_PARSE
    end
    wire [ARBT_NUM-1:0] burst_mask_nxt;
    wire burst_mask_ena;
    wire burst_mask_set;
    wire burst_mask_clr;
      assign burst_mask_set = o_icb_cmd_beat[0] & arbt_ena;
      assign burst_mask_clr = (|burst_mask_r) & o_icb_cmd_beat[1] & arbt_ena;
    assign burst_mask_ena = clk_en & (burst_mask_set | burst_mask_clr);
    assign burst_mask_nxt = burst_mask_clr ? {ARBT_NUM{1'b0}} : (~i_bus_icb_cmd_sel); 
e603_subsys_gnrl_dfflr #(ARBT_NUM) burst_mask_dfflr (burst_mask_ena, burst_mask_nxt, burst_mask_r, clk, rst_n);// VPP_NO_REG_PARSE
      assign i_bus_icb_cmd_valid_pos   = (~burst_mask_r) & (~omask_r) & (~lock_mask_r) & i_bus_icb_cmd_valid;
      assign i_bus_icb_cmd_ready       = (~burst_mask_r) & (~omask_r) & (~lock_mask_r) & i_bus_icb_cmd_ready_pos;
      assign i_bus_icb_cmd_sel_vec_pos = (~burst_mask_r) & (~omask_r) & (~lock_mask_r) & i_bus_icb_cmd_sel_vec;
    assign o_icb_cmd_sel   = |i_bus_icb_cmd_sel_vec_pos;
    assign o_icb_cmd_valid = o_icb_cmd_valid_real & (~rspid_fifo_full);
    assign o_icb_cmd_ready_real = o_icb_cmd_ready & (~rspid_fifo_full);
    for(i = 0; i < ARBT_NUM; i = i+1)
    begin:gen_icb_distract
      assign i_icb_cmd_read [i] = i_bus_icb_cmd_read [(i+1)*1     -1 : i*1     ];
      assign i_icb_cmd_addr [i] = i_bus_icb_cmd_addr [(i+1)*AW    -1 : i*AW    ];
      assign i_icb_cmd_wdata[i] = i_bus_icb_cmd_wdata[(i+1)*DW    -1 : i*DW    ];
      assign i_icb_cmd_wmask[i] = i_bus_icb_cmd_wmask[(i+1)*DW/8    -1 : i*DW/8    ];
      assign i_icb_cmd_beat [i] = i_bus_icb_cmd_beat [(i+1)*2     -1 : i*2     ];
      assign i_icb_cmd_lock [i] = i_bus_icb_cmd_lock [(i+1)*1     -1 : i*1     ];
      assign i_icb_cmd_excl [i] = i_bus_icb_cmd_excl [(i+1)*1     -1 : i*1     ];
      assign i_icb_cmd_size [i] = i_bus_icb_cmd_size [(i+1)*CMD_SIZE_W     -1 : i*CMD_SIZE_W     ];
      assign i_icb_cmd_usr  [i] = i_bus_icb_cmd_usr  [(i+1)*CMD_UW -1 : i*CMD_UW ];
      assign i_icb_cmd_id   [i] = i_bus_icb_cmd_id   [(i+1)*ID_W -1 : i*ID_W ];
      assign i_icb_cmd_xlen  [i] = i_bus_icb_cmd_xlen   [(i+1)*8 -1 : i*8 ];
      assign i_icb_cmd_xburst[i] = i_bus_icb_cmd_xburst [(i+1)*2 -1 : i*2 ];
      assign i_icb_cmd_modes [i] = i_bus_icb_cmd_modes  [(i+1)*2 -1 : i*2 ];
      assign i_icb_cmd_dmode [i] = i_bus_icb_cmd_dmode  [(i+1)*1 -1 : i*1 ];
      assign i_icb_cmd_attri [i] = i_bus_icb_cmd_attri  [(i+1)*3 -1 : i*3 ];
      assign i_bus_icb_cmd_ready_pos[i] = i_bus_icb_cmd_grt_vec[i] & o_icb_cmd_ready_real;
      assign i_bus_icb_rsp_valid[i] = icb_rsp_valid_pre & (icb_rsp_port_id == i[ARBT_PTR_W-1:0]);
    end
    assign arbt_ena = o_icb_cmd_valid & o_icb_cmd_ready;
      wire [ARBT_NUM-1:0] lock_mask_set;
      wire [ARBT_NUM-1:0] lock_mask_clr;
      wire [ARBT_NUM-1:0] lock_mask_ena;
      wire [ARBT_NUM-1:0] lock_mask_nxt;
      for(i = 0; i < ARBT_NUM; i = i+1) begin:gen_lock_mask
        assign lock_mask_set[i] = clk_en & (i_bus_icb_cmd_sel[i] == 1'b0) & o_icb_cmd_lock & arbt_ena;
        assign lock_mask_clr[i] = clk_en & lock_mask_r[i] & ((~o_icb_cmd_lock) & arbt_ena);
        assign lock_mask_ena[i] = lock_mask_set[i] |   lock_mask_clr[i];
        assign lock_mask_nxt[i] = lock_mask_set[i] & (~lock_mask_clr[i]);
        if(SUPPORT_LOCK == 1) begin: support_lock_gen
e603_subsys_gnrl_dfflr #(1) lock_mask_dfflr (lock_mask_ena[i], lock_mask_nxt[i], lock_mask_r[i], clk, rst_n);// VPP_NO_REG_PARSE
        end
        else begin: no_support_lock_gen
        assign lock_mask_r[i] = 1'b0;
        end
      end
    if(ARBT_SCHEME == ARBT_SCHEME_PRIORITY) begin:gen_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_icb_cmd_grt_vec[i] =  1'b1;
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_valid_pos[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_icb_cmd_grt_vec[i] =  ~(|i_bus_icb_cmd_valid_pos[i-1:0]);
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_valid_pos[i];
        end
      end
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN) begin:gen_rrobin_arbt
       if(RRBIN_CUT_TIMING == 1) begin:gen_rbin_cut_timing
      wire lock_mask_r_set  = |(lock_mask_set & (~lock_mask_clr));
      wire burst_mask_r_set = |(burst_mask_set & (~burst_mask_clr));
     e603_subsys_gnrl_rrobin_cut # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin_cut(
       .rrobin_active (rrobin_notime_active),
       .grt_vec  (i_bus_icb_cmd_grt_vec),
       .req_vec  (i_bus_icb_cmd_sel_vec_pos),
       .req_mask  (burst_mask_r | lock_mask_r),
       .req_mask_set  (burst_mask_r_set | lock_mask_r_set),
       .arbt_ena (arbt_ena & clk_en),
       .clk      (clk),
       .rst_n    (rst_n)
     );
       end
       else begin: no_gen_rbin_cut_ciming
     e603_subsys_gnrl_rrobin # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin(
       .rrobin_active (rrobin_notime_active),
       .grt_vec  (i_bus_icb_cmd_grt_vec),
       .req_vec  (i_bus_icb_cmd_sel_vec_pos),
       .arbt_ena (arbt_ena & clk_en),
       .clk      (clk),
       .rst_n    (rst_n)
     );
       end
     assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec;
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
   end
   else begin: gen_no_rrobin
     assign rrobin_notime_active = 1'b0;
   end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN_TIME) begin:gen_rrobin_time_arbt
     e603_subsys_gnrl_rrobin_time # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin_time(
       .rrobin_active (rrobin_time_active),
       .grt_vec  (i_bus_icb_cmd_grt_vec),
       .req_vec  (i_bus_icb_cmd_valid),
       .req_mask  (burst_mask_r | lock_mask_r),
       .arbt_ena (arbt_ena & clk_en),
       .clk      (clk),
       .rst_n    (rst_n)
     );
     assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec;
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid & i_bus_icb_cmd_sel);
   end
   else begin: gen_no_rrobin_time
     assign rrobin_time_active = 1'b0;
   end
   assign rrobin_active = rrobin_notime_active | rrobin_time_active | rbin4_active;
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_1HOT) begin:gen_indic_arbt
     assign i_bus_icb_cmd_grt_vec = i_bus_icb_cmd_sel_vec_pos;
     assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec;
     assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
   end
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_PRIORITY) begin:gen_indic_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_icb_cmd_grt_vec[i] =  1'b1;
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_sel_vec_pos[i];
        end
        else if(i==(ARBT_NUM-1)) begin: gen_i_is_n
          assign i_bus_icb_cmd_grt_vec[i] =  ~(|i_bus_icb_cmd_sel_vec_pos[i-1:0]);
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_icb_cmd_grt_vec[i] =  ~(|i_bus_icb_cmd_sel_vec_pos[i-1:0]);
          assign i_bus_icb_cmd_sel[i] = i_bus_icb_cmd_grt_vec[i] & i_bus_icb_cmd_sel_vec_pos[i];
        end
      end
      assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN4) begin:gen_rbin4_arbt
      wire lock_mask_r_set  = |lock_mask_set ;
      wire burst_mask_r_set = |burst_mask_set;
      e603_subsys_gnrl_rbin4 # (
          .ARBT_NUM(ARBT_NUM)
      )u_e603_subsys_gnrl_rbin4(
        .grt_vec  (i_bus_icb_cmd_grt_vec),
        .req_vec  (i_bus_icb_cmd_sel_vec_pos),
        .arbt_ena (arbt_ena & clk_en & (~lock_mask_r_set) & (~burst_mask_r_set)),
        .rbin4_active(rbin4_active),
        .clk      (clk),
        .rst_n    (rst_n)
      );
      assign i_bus_icb_cmd_sel = i_bus_icb_cmd_grt_vec & i_bus_icb_cmd_sel_vec_pos;
      assign o_icb_cmd_valid_real = |(i_bus_icb_cmd_valid_pos & i_bus_icb_cmd_sel);
   end
   else begin:gen_no_rbin4_arbt
      assign rbin4_active = 1'b0;
   end
    always @ (*) begin : sel_o_icb_cmd_ready_PROC
      sel_o_icb_cmd_read  = {1   {1'b0}};
      sel_o_icb_cmd_addr  = {AW  {1'b0}};
      sel_o_icb_cmd_wdata = {DW  {1'b0}};
      sel_o_icb_cmd_wmask = {DW/8  {1'b0}};
      sel_o_icb_cmd_beat  = {2   {1'b0}};
      sel_o_icb_cmd_lock  = {1   {1'b0}};
      sel_o_icb_cmd_excl  = {1   {1'b0}};
      sel_o_icb_cmd_size  = {CMD_SIZE_W   {1'b0}};
      sel_o_icb_cmd_usr   = {CMD_UW{1'b0}};
      sel_o_icb_cmd_id    = {ID_W{1'b0}};
      sel_o_icb_cmd_xlen  = {8{1'b0}};
      sel_o_icb_cmd_xburst= {2{1'b0}};
      sel_o_icb_cmd_modes = {2{1'b0}};
      sel_o_icb_cmd_dmode = {1{1'b0}};
      sel_o_icb_cmd_attri = {3{1'b0}};
      for(j = 0; j < ARBT_NUM; j = j+1) begin
        sel_o_icb_cmd_read  = sel_o_icb_cmd_read  | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_read [j]);
        sel_o_icb_cmd_addr  = sel_o_icb_cmd_addr  | ({AW   {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_addr [j]);
        sel_o_icb_cmd_wdata = sel_o_icb_cmd_wdata | ({DW   {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_wdata[j]);
        sel_o_icb_cmd_wmask = sel_o_icb_cmd_wmask | ({DW/8   {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_wmask[j]);
        sel_o_icb_cmd_beat  = sel_o_icb_cmd_beat  | ({2    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_beat [j]);
        sel_o_icb_cmd_lock  = sel_o_icb_cmd_lock  | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_lock [j]);
        sel_o_icb_cmd_excl  = sel_o_icb_cmd_excl  | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_excl [j]);
        sel_o_icb_cmd_size  = sel_o_icb_cmd_size  | ({CMD_SIZE_W    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_size [j]);
        sel_o_icb_cmd_usr   = sel_o_icb_cmd_usr   | ({CMD_UW{i_bus_icb_cmd_sel[j]}} & i_icb_cmd_usr  [j]);
        sel_o_icb_cmd_id    = sel_o_icb_cmd_id    | ({ID_W  {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_id   [j]);
        sel_o_icb_cmd_xlen  = sel_o_icb_cmd_xlen  | ({8    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_xlen  [j]);
        sel_o_icb_cmd_xburst= sel_o_icb_cmd_xburst| ({2    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_xburst[j]);
        sel_o_icb_cmd_modes = sel_o_icb_cmd_modes | ({2    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_modes [j]);
        sel_o_icb_cmd_dmode = sel_o_icb_cmd_dmode | ({1    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_dmode [j]);
        sel_o_icb_cmd_attri = sel_o_icb_cmd_attri | ({3    {i_bus_icb_cmd_sel[j]}} & i_icb_cmd_attri [j]);
      end
    end
    always @ (*) begin : i_arbt_indic_id_PROC
      i_arbt_indic_id = {ARBT_PTR_W{1'b0}};
      for(j = 0; j < ARBT_NUM; j = j+1) begin
// spyglass disable_block W216
// SMD: Inappropriate range select for int_part_sel variable
// SJ:  Here is not a real issue
        i_arbt_indic_id = i_arbt_indic_id | ({ARBT_PTR_W{i_bus_icb_cmd_sel[j]}} & (j[ARBT_PTR_W-1:0]));
// spyglass enable_block W216
      end
    end
    assign rspid_fifo_wen = 1'b0;
    assign rspid_fifo_ren = 1'b0;
    if(ALLOW_0CYCL_RSP == 1) begin: gen_allow_0rsp
        assign rspid_fifo_bypass = rspid_fifo_empty & rspid_fifo_wen & rspid_fifo_ren;
        if(I_ICB_IDW_ZERO == 1) begin: rsp_port_id_i_idw0
            assign icb_rsp_port_id = rspid_fifo_empty ? rspid_fifo_wdat : icb_rsp_id;
        end
        else begin: rsp_port_id_i_idwx
            if(I_REAL_ID_W != 0) begin: rsp_port_id_i_idw_not0
                assign icb_rsp_port_id = rspid_fifo_empty ? rspid_fifo_wdat : icb_rsp_id[I_REAL_ID_W+ARBT_PTR_W-1:I_REAL_ID_W];
            end
            else begin: rsp_port_id_i_idw_is0
                assign icb_rsp_port_id = rspid_fifo_empty ? rspid_fifo_wdat : icb_rsp_id[ID_W-1:ID_W-ARBT_PTR_W];
            end
        end
        assign icb_rsp_valid_pre = icb_rsp_valid;
        assign icb_rsp_ready     = icb_rsp_ready_pre;
    end
    else begin: gen_no_allow_0rsp
        assign rspid_fifo_bypass   = 1'b0;
        if(I_ICB_IDW_ZERO == 1) begin: rsp_port_id_i_idw0
            assign icb_rsp_port_id   = icb_rsp_id;
        end
        else begin: rsp_port_id_i_idwx
            if(I_REAL_ID_W != 0) begin: rsp_port_id_i_idw_not0
                assign icb_rsp_port_id   = icb_rsp_id[I_REAL_ID_W+ARBT_PTR_W-1:I_REAL_ID_W];
            end
            else begin: rsp_port_id_i_idw_is0
                assign icb_rsp_port_id   = icb_rsp_id[ID_W-1:ID_W-ARBT_PTR_W];
            end
        end
        assign icb_rsp_valid_pre = icb_rsp_valid;
        assign icb_rsp_ready     = icb_rsp_ready_pre;
    end
    assign rspid_fifo_i_valid = clk_en & rspid_fifo_wen & (~rspid_fifo_bypass);
    assign rspid_fifo_full    = (~rspid_fifo_i_ready);
    assign rspid_fifo_o_ready = clk_en & rspid_fifo_ren & (~rspid_fifo_bypass);
    assign rspid_fifo_empty   = (~rspid_fifo_o_valid);
    assign rspid_fifo_wdat   = i_arbt_indic_id;
    if(FIFO_OUTS_NUM == 1) begin:gen_dp_1
      e603_subsys_gnrl_pipe_stage # (
        .CUT_READY (FIFO_CUT_READY),
        .DP  (1),
        .DW  (ARBT_PTR_W)
      ) u_e603_subsys_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else begin: gen_dp_gt1
      e603_subsys_gnrl_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT(FIFO_REG_OUT),
        .CUT_READY(FIFO_CUT_READY),
        .DP  (FIFO_OUTS_NUM),
        .DW  (ARBT_PTR_W)
      ) u_e603_subsys_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    assign o_icb_cmd_read  = sel_o_icb_cmd_read ;
    assign o_icb_cmd_addr  = sel_o_icb_cmd_addr ;
    assign o_icb_cmd_wdata = sel_o_icb_cmd_wdata;
    assign o_icb_cmd_wmask = sel_o_icb_cmd_wmask;
    assign o_icb_cmd_beat  = sel_o_icb_cmd_beat ;
    assign o_icb_cmd_lock  = sel_o_icb_cmd_lock ;
    assign o_icb_cmd_excl  = sel_o_icb_cmd_excl ;
    assign o_icb_cmd_size  = sel_o_icb_cmd_size ;
    assign o_icb_cmd_usr   = sel_o_icb_cmd_usr  ;
        if(I_ICB_IDW_ZERO == 1) begin: cmd_id_i_idw0
    assign o_icb_cmd_id    = rspid_fifo_wdat[ARBT_PTR_W-1:0];
        end
        else begin: cmd_id_i_idwx
            if(I_REAL_ID_W != 0) begin: cmd_id_id_i_idw_not0
                  if((ARBT_PTR_W+I_REAL_ID_W) < ID_W) begin: ptr_w_rlidw_lt_idw
    assign o_icb_cmd_id    = {{ID_W-ARBT_PTR_W-I_REAL_ID_W{1'b0}},
                              rspid_fifo_wdat[ARBT_PTR_W-1:0], sel_o_icb_cmd_id[I_REAL_ID_W-1:0]};
                  end
                  else begin: ptr_w_rlidw_eq_idw
    assign o_icb_cmd_id    = {rspid_fifo_wdat[ARBT_PTR_W-1:0], sel_o_icb_cmd_id[I_REAL_ID_W-1:0]};
                  end
            end
            else begin: cmd_id_id_i_idw_is0
    assign o_icb_cmd_id    = {rspid_fifo_wdat[ARBT_PTR_W-1:0], sel_o_icb_cmd_id[ID_W-ARBT_PTR_W-1:0]};
            end
        end
    assign o_icb_cmd_xlen  = sel_o_icb_cmd_xlen  ;
    assign o_icb_cmd_xburst= sel_o_icb_cmd_xburst;
    assign o_icb_cmd_modes = sel_o_icb_cmd_modes ;
    assign o_icb_cmd_dmode = sel_o_icb_cmd_dmode ;
    assign o_icb_cmd_attri = sel_o_icb_cmd_attri ;
    assign icb_rsp_ready_pre = i_bus_icb_rsp_ready[icb_rsp_port_id];
    assign i_bus_icb_rsp_err     = {ARBT_NUM{icb_rsp_err  }};
    assign i_bus_icb_rsp_excl_ok = {ARBT_NUM{icb_rsp_excl_ok}};
    assign i_bus_icb_rsp_rdata   = {ARBT_NUM{icb_rsp_rdata}};
    assign i_bus_icb_rsp_usr     = {ARBT_NUM{icb_rsp_usr}};
    wire[ID_W-1:0] icb_rsp_id_ext;
        if(I_ICB_IDW_ZERO == 1) begin: rsp_id_i_idw0
    assign icb_rsp_id_ext = {ID_W{1'b0}};
        end
        else begin: rsp_id_i_idwx
            if(I_REAL_ID_W != 0) begin: rsp_id_i_idw_not0
    assign icb_rsp_id_ext = { {ID_W-I_REAL_ID_W{1'b0}}, icb_rsp_id[I_REAL_ID_W-1:0] };
            end
            else begin: rsp_id_i_idw_is0
    assign icb_rsp_id_ext = { {ARBT_PTR_W{1'b0}}, icb_rsp_id[ID_W-ARBT_PTR_W-1:0] };
            end
        end
    assign i_bus_icb_rsp_id      = {ARBT_NUM{ icb_rsp_id_ext }};
    assign i_bus_icb_rsp_last    = {ARBT_NUM{icb_rsp_last}};
  end
  endgenerate 
  assign arbt_active =
         (|i_bus_icb_cmd_sel_vec) | (~rspid_fifo_empty) | icb_rsp_valid | (|burst_mask_r)| (|omask_r) | (|lock_mask_r) | rrobin_active;
endmodule
module e603_subsys_gnrl_ficb_buffer_id # (
    parameter OUTS_CNT_BLOCK_THROUGH = 0,
    parameter ID_W = 4,
    parameter RSP_STRICT_ORDER = 1,
  parameter PAYLOAD_NORST = 0,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter CMD_MSKO = 0,
  parameter OUTS_CNT_W = 1,
  parameter AW = 32,
  parameter DW = 32,
  parameter CMD_CUT_READY = 0,
  parameter RSP_CUT_READY = 0,
  parameter ACTIVE_USE_FLOP_CLEAN = 0,
  parameter CMD_DP = 0,
  parameter RSP_DP = 0,
  parameter CMD_BYPBUF = 0,
  parameter CMD_RGLR_FIFO = 0,
  parameter RSP_BYPBUF = 0,
  parameter RSP_RGLR_FIFO = 0,
  parameter REG_OUT = 0,
  parameter RSP_ALWAYS_READY = 0,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  input              i_clk_en,
  input              o_clk_en,
  output             icb_buffer_active,
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [DW-1:0]    i_icb_cmd_wdata,
  input  [DW/8-1:0]  i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  input  [ID_W-1:0] i_icb_cmd_id,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [DW-1:0]    i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [DW-1:0]    o_icb_cmd_wdata,
  output [DW/8-1:0]  o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  output [ID_W-1:0] o_icb_cmd_id,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  localparam CMD_PACK_W = (1+AW+DW+DW/8+1+3+3+CMD_UW+8+2+2+1+3+ID_W + 0);
  localparam RSP_PACK_W = (2+DW+RSP_UW+ID_W+1 + 0);
 wire i_icb_cmd_xlen_eq0 = (i_icb_cmd_xlen == 8'd0);
 wire i_icb_cmd_first = i_icb_cmd_beat[0] | i_icb_cmd_xlen_eq0;
 wire o_icb_cmd_xlen_eq0 = (o_icb_cmd_xlen == 8'd0);
 wire o_icb_cmd_first = o_icb_cmd_beat[0] | o_icb_cmd_xlen_eq0;
 generate
   if((CMD_DP == 0) && (RSP_DP == 0)) begin:gen_icb_buf_through
  wire outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready & i_clk_en 
    ;
  wire outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & i_clk_en 
    ;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
      assign icb_buffer_active =
      i_icb_cmd_sel | (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
    wire i_outs_cnt_is_max;
    if(OUTS_CNT_BLOCK_THROUGH == 1) begin:outs_cnt_block_through
        assign i_outs_cnt_is_max = (outs_cnt_r == {OUTS_CNT_W{1'b1}});
    end
    else begin:outs_cnt_no_block_through
        assign i_outs_cnt_is_max = 1'b0;
    end
    assign i_icb_cmd_ready = (~i_outs_cnt_is_max) & o_icb_cmd_ready;
    assign o_icb_cmd_sel   = (~i_outs_cnt_is_max) & i_icb_cmd_sel;
    assign o_icb_cmd_valid = (~i_outs_cnt_is_max) & i_icb_cmd_valid;
    assign o_icb_cmd_read  = i_icb_cmd_read ;
    assign o_icb_cmd_addr  = i_icb_cmd_addr ;
    assign o_icb_cmd_wdata = i_icb_cmd_wdata;
    assign o_icb_cmd_wmask = i_icb_cmd_wmask;
    assign o_icb_cmd_beat  = i_icb_cmd_beat ;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
    assign o_icb_cmd_size  = o_icb_cmd_size_pre ;
    assign o_icb_cmd_xlen  = o_icb_cmd_xlen_pre  ;
    assign o_icb_cmd_lock  = i_icb_cmd_lock ;
    assign o_icb_cmd_excl  = i_icb_cmd_excl ;
    assign o_icb_cmd_size_pre  = i_icb_cmd_size ;
    assign o_icb_cmd_usr   = i_icb_cmd_usr  ;
    assign o_icb_cmd_id    = i_icb_cmd_id  ;
    assign o_icb_cmd_xlen_pre  = i_icb_cmd_xlen  ;
    assign o_icb_cmd_xburst= i_icb_cmd_xburst;
    assign o_icb_cmd_modes = i_icb_cmd_modes ;
    assign o_icb_cmd_dmode = i_icb_cmd_dmode ;
    assign o_icb_cmd_attri = i_icb_cmd_attri ;
    assign o_icb_rsp_ready = i_icb_rsp_ready;
    assign i_icb_rsp_valid     = o_icb_rsp_valid;
    assign i_icb_rsp_err       = o_icb_rsp_err  ;
    assign i_icb_rsp_excl_ok   = o_icb_rsp_excl_ok  ;
    assign i_icb_rsp_rdata     = o_icb_rsp_rdata;
    assign i_icb_rsp_usr       = o_icb_rsp_usr;
    assign i_icb_rsp_id        = o_icb_rsp_id ;
    assign i_icb_rsp_last        = o_icb_rsp_last ;
  end
  else begin:gen_icb_buf_not_through
  wire [CMD_PACK_W-1:0] cmd_fifo_i_dat = {
                                 i_icb_cmd_read,
                                 i_icb_cmd_addr,
                                 i_icb_cmd_wdata,
                                 i_icb_cmd_wmask,
                                 i_icb_cmd_lock,
                                 i_icb_cmd_excl,
                                 i_icb_cmd_size,
                                 i_icb_cmd_beat,
                                 i_icb_cmd_xlen,
                                 i_icb_cmd_xburst,
                                 i_icb_cmd_modes,
                                 i_icb_cmd_dmode,
                                 i_icb_cmd_attri,
                                 i_icb_cmd_id,
                                 i_icb_cmd_usr};
  wire [CMD_PACK_W-1:0] cmd_fifo_o_dat;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
    assign o_icb_cmd_size  = o_icb_cmd_size_pre ;
    assign o_icb_cmd_xlen  = o_icb_cmd_xlen_pre  ;
  assign {
                                 o_icb_cmd_read,
                                 o_icb_cmd_addr,
                                 o_icb_cmd_wdata,
                                 o_icb_cmd_wmask,
                                 o_icb_cmd_lock,
                                 o_icb_cmd_excl,
                                 o_icb_cmd_size_pre,
                                 o_icb_cmd_beat,
                                 o_icb_cmd_xlen_pre,
                                 o_icb_cmd_xburst,
                                 o_icb_cmd_modes,
                                 o_icb_cmd_dmode,
                                 o_icb_cmd_attri,
                                 o_icb_cmd_id,
                                 o_icb_cmd_usr} = cmd_fifo_o_dat;
  wire o_icb_cmd_valid_pre;
  wire o_icb_cmd_ready_pre;
  wire outs_cnt_full;
  wire cmd_fifo_i_valid;
  wire cmd_fifo_i_ready;
  assign cmd_fifo_i_valid = (~outs_cnt_full) & i_icb_cmd_valid;
  assign i_icb_cmd_ready  = (~outs_cnt_full) & cmd_fifo_i_ready;
  wire cmd_ratio_fifo_active;
    if(CMD_RGLR_FIFO == 1) begin: gen_cmd_rlgr_fifo
  e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP  (CMD_DP),
    .DW  (CMD_PACK_W)
  ) u_e603_subsys_gnrl_cmd_fifo (
    .i_vld(cmd_fifo_i_valid),
    .i_rdy(cmd_fifo_i_ready),
    .i_dat(cmd_fifo_i_dat ),
    .o_vld(o_icb_cmd_valid_pre),
    .o_rdy(o_icb_cmd_ready_pre),
    .o_dat(cmd_fifo_o_dat ),
    .clk  (clk),
    .rst_n(rst_n)
  );
   assign cmd_ratio_fifo_active = o_icb_cmd_valid_pre;
    end
    else if(CMD_BYPBUF == 0) begin: gen_cmd_no_bypbuf
  e603_subsys_gnrl_ratio_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .I_SUPPORT_RATIO (I_SUPPORT_RATIO),
        .O_SUPPORT_RATIO (O_SUPPORT_RATIO),
    .DP  (CMD_DP),
    .DW  (CMD_PACK_W)
  ) u_e603_subsys_gnrl_cmd_fifo (
    .i_clk_en     (i_clk_en),
    .o_clk_en     (o_clk_en),
    .o_fifo_active(cmd_ratio_fifo_active),
    .i_vld(cmd_fifo_i_valid),
    .i_rdy(cmd_fifo_i_ready),
    .i_dat(cmd_fifo_i_dat ),
    .o_vld(o_icb_cmd_valid_pre),
    .o_rdy(o_icb_cmd_ready_pre),
    .o_dat(cmd_fifo_o_dat ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    else begin:gen_cmd_bypbuf
  e603_subsys_gnrl_bypbuf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP  (CMD_DP),
    .DW  (CMD_PACK_W)
  ) u_e603_subsys_gnrl_cmd_bypbuf (
    .i_vld(cmd_fifo_i_valid & i_clk_en),
    .i_rdy(cmd_fifo_i_ready),
    .i_dat(cmd_fifo_i_dat ),
    .o_vld(o_icb_cmd_valid_pre),
    .o_rdy(o_icb_cmd_ready_pre & o_clk_en),
    .o_dat(cmd_fifo_o_dat ),
        .fifo_o_vld(cmd_ratio_fifo_active),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
   wire oo_outs_cnt_max;
   wire o_outs_cnt_max;
    if(CMD_DP == 0) begin:dp_is_0_gen
        assign o_icb_cmd_sel = i_icb_cmd_sel;
    end
    else begin:dp_is_not_0_gen
        assign o_icb_cmd_sel = o_icb_cmd_valid_pre;
    end
  wire rsp_buf_ready;
    if(RSP_ALWAYS_READY == 1) begin: gen_rsp_always_ready_1
      assign o_icb_cmd_valid     = rsp_buf_ready & o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = rsp_buf_ready & o_icb_cmd_ready;
    end
    else begin: gen_rsp_always_ready_0
      assign o_icb_cmd_valid     = o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = o_icb_cmd_ready;
    end
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata,
                                 o_icb_rsp_id,
                                 o_icb_rsp_last,
                                 o_icb_rsp_usr};
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 i_icb_rsp_err,
                                 i_icb_rsp_excl_ok,
                                 i_icb_rsp_rdata,
                                 i_icb_rsp_id,
                                 i_icb_rsp_last,
                                 i_icb_rsp_usr} = rsp_fifo_o_dat;
  wire o_icb_rsp_valid_raw;
  wire o_icb_rsp_ready_raw;
    if(RSP_RGLR_FIFO == 1) begin: gen_rsp_rlgr_fifo
      e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT (REG_OUT),
        .DP  (RSP_DP),
        .DW  (RSP_PACK_W)
      ) u_e603_subsys_gnrl_rsp_fifo (
        .i_vld(o_icb_rsp_valid_raw),
        .i_rdy(o_icb_rsp_ready_raw),
        .i_dat(rsp_fifo_i_dat ),
        .o_vld(i_icb_rsp_valid),
        .o_rdy(i_icb_rsp_ready),
        .o_dat(rsp_fifo_o_dat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else if(RSP_BYPBUF == 0) begin: gen_rsp_no_bypbuf
      e603_subsys_gnrl_ratio_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .I_SUPPORT_RATIO (O_SUPPORT_RATIO),
        .O_SUPPORT_RATIO (I_SUPPORT_RATIO),
        .REG_OUT (REG_OUT),
        .DP  (RSP_DP),
        .DW  (RSP_PACK_W)
      ) u_e603_subsys_gnrl_rsp_fifo (
        .i_clk_en     (o_clk_en),
        .o_clk_en     (i_clk_en),
        .o_fifo_active(),
        .i_vld(o_icb_rsp_valid_raw),
        .i_rdy(o_icb_rsp_ready_raw),
        .i_dat(rsp_fifo_i_dat ),
        .o_vld(i_icb_rsp_valid),
        .o_rdy(i_icb_rsp_ready),
        .o_dat(rsp_fifo_o_dat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else begin:gen_rsp_bypbuf
      e603_subsys_gnrl_bypbuf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RSP_DP),
        .DW  (RSP_PACK_W)
      ) u_e603_subsys_gnrl_rsp_bypbuf (
        .i_vld(o_icb_rsp_valid_raw & o_clk_en),
        .i_rdy(o_icb_rsp_ready_raw),
        .i_dat(rsp_fifo_i_dat ),
        .o_vld(i_icb_rsp_valid),
        .o_rdy(i_icb_rsp_ready & i_clk_en),
        .o_dat(rsp_fifo_o_dat ),
        .fifo_o_vld(),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
  wire outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready & i_clk_en
                    ;
  wire outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & i_clk_en
                    ;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign outs_cnt_full = (outs_cnt_r == {OUTS_CNT_W{1'b1}});
   if((CMD_BYPBUF != 1) && (CMD_DP != 0) && (ACTIVE_USE_FLOP_CLEAN == 1)) begin:gen_active_flop_clean
  assign icb_buffer_active =
      (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
   end
   else begin: gen_active_no_flop_clean
  assign icb_buffer_active =
      i_icb_cmd_sel | cmd_ratio_fifo_active | (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
   end
  wire o_outs_cnt_inc = o_icb_cmd_valid & o_icb_cmd_ready & o_clk_en 
                    ;
  wire o_outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & i_clk_en 
                    ;
  wire o_outs_cnt_ena = o_outs_cnt_inc ^ o_outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_r;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_nxt = o_outs_cnt_inc ? (o_outs_cnt_r + 1'b1) : (o_outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) o_outs_cnt_dfflr (o_outs_cnt_ena, o_outs_cnt_nxt, o_outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire [OUTS_CNT_W-1:0] o_outs_cnt_din = o_outs_cnt_ena ? o_outs_cnt_nxt : o_outs_cnt_r;
  wire rsp_buf_ready_raw = ~(o_outs_cnt_r   == RSP_DP[OUTS_CNT_W-1:0]);
  wire rsp_buf_ready_din = ~(o_outs_cnt_din == RSP_DP[OUTS_CNT_W-1:0]);
    wire o_need_updat = o_outs_cnt_ena;
    wire o_need_updat_r;
    wire o_need_updat_r_set = (o_need_updat && !o_clk_en);
    wire o_need_updat_r_clr = (o_need_updat_r && o_clk_en);
    wire o_need_updat_r_ena = o_need_updat_r_set || o_need_updat_r_clr;
    wire o_need_updat_r_nxt = o_need_updat_r_set;
e603_subsys_gnrl_dfflr  #(1) o_need_updat_r_dfflr    (o_need_updat_r_ena, o_need_updat_r_nxt, o_need_updat_r,     clk, rst_n);// VPP_NO_REG_PARSE
    wire rsp_buf_ready_r;
    wire rsp_buf_ready_r_ena = o_clk_en && (o_need_updat || o_need_updat_r);
    wire rsp_buf_ready_r_nxt = (o_need_updat ? rsp_buf_ready_din : rsp_buf_ready_raw);
e603_subsys_gnrl_dfflrs  #(1) rsp_buf_ready_r_dfflrs    (rsp_buf_ready_r_ena, rsp_buf_ready_r_nxt, rsp_buf_ready_r,     clk, rst_n);// VPP_NO_REG_PARSE
  assign rsp_buf_ready = rsp_buf_ready_r;
  wire oo_outs_cnt_inc = o_icb_cmd_valid & o_icb_cmd_ready & o_clk_en 
                    ;
  wire oo_outs_cnt_dec = o_icb_rsp_valid & o_icb_rsp_ready & o_clk_en 
                    ;
  wire oo_outs_cnt_ena = oo_outs_cnt_inc ^ oo_outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] oo_outs_cnt_r;
  wire [OUTS_CNT_W-1:0] oo_outs_cnt_nxt = oo_outs_cnt_inc ? (oo_outs_cnt_r + 1'b1) : (oo_outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) oo_outs_cnt_dfflr (oo_outs_cnt_ena, oo_outs_cnt_nxt, oo_outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire oo_outs_cnt_eq0 = (oo_outs_cnt_r == {OUTS_CNT_W{1'b0}});
  assign oo_outs_cnt_max = (oo_outs_cnt_r == {OUTS_CNT_W{1'b1}});
  assign o_outs_cnt_max = (o_outs_cnt_r == {OUTS_CNT_W{1'b1}});
  if (RSP_STRICT_ORDER == 1) begin: rsp_strict_order_gen
      assign o_icb_rsp_valid_raw = (~oo_outs_cnt_eq0) & o_icb_rsp_valid;
      assign o_icb_rsp_ready     = (~oo_outs_cnt_eq0) & o_icb_rsp_ready_raw;
  end
  else begin: rsp_no_order_gen
      assign o_icb_rsp_valid_raw = o_icb_rsp_valid;
      assign o_icb_rsp_ready     = o_icb_rsp_ready_raw;
  end
  end
  endgenerate
endmodule
module e603_subsys_gnrl_ficb_async_id # (
    parameter ID_W = 4,
    parameter RSP_STRICT_ORDER = 1,
  parameter PAYLOAD_NORST = 0,
  parameter RSP_ALWAYS_READY = 0,
  parameter OUTS_CNT_W = 1,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 4,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter AW = 32,
  parameter DW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  output             icb2icb_async_i_active,
  output             icb2icb_async_o_active,
  input              i_icb_cmd_sel  ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [DW-1:0]    i_icb_cmd_wdata,
  input  [DW/8-1:0]    i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [ID_W-1:0] i_icb_cmd_id,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [DW-1:0]    i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel  ,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [DW-1:0]    o_icb_cmd_wdata,
  output [DW/8-1:0]    o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input              i_clk,
  input              o_clk,
  input              i_rst_n,
  input              o_rst_n
  );
 wire i_icb_cmd_xlen_eq0 = (i_icb_cmd_xlen == 8'd0);
 wire i_icb_cmd_first = i_icb_cmd_beat[0] | i_icb_cmd_xlen_eq0;
 wire o_icb_cmd_xlen_eq0 = (o_icb_cmd_xlen == 8'd0);
 wire o_icb_cmd_first = o_icb_cmd_beat[0] | o_icb_cmd_xlen_eq0;
  wire i_icb_reset_flag_r;
e603_subsys_gnrl_dffrs #(1) reset_flag_dffrs (1'b0, i_icb_reset_flag_r, i_clk, i_rst_n);// VPP_NO_REG_PARSE
  localparam CMD_PACK_W = (1+AW+DW+DW/8+1+4+2+CMD_UW+8+2+2+1+3+ID_W+0);
  wire [CMD_PACK_W-1:0] cmd_fifo_i_dat = {
                                 i_icb_cmd_read,
                                 i_icb_cmd_addr,
                                 i_icb_cmd_wdata,
                                 i_icb_cmd_wmask,
                                 i_icb_cmd_lock,
                                 i_icb_cmd_excl,
                                 i_icb_cmd_size,
                                 i_icb_cmd_beat,
                                 i_icb_cmd_xlen,
                                 i_icb_cmd_xburst,
                                 i_icb_cmd_modes,
                                 i_icb_cmd_dmode,
                                 i_icb_cmd_attri,
                                 i_icb_cmd_id,
                                 i_icb_cmd_usr};
  wire [CMD_PACK_W-1:0] cmd_fifo_o_dat;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
    assign o_icb_cmd_size  = o_icb_cmd_size_pre ;
    assign o_icb_cmd_xlen  = o_icb_cmd_xlen_pre  ;
  assign {
                                 o_icb_cmd_read,
                                 o_icb_cmd_addr,
                                 o_icb_cmd_wdata,
                                 o_icb_cmd_wmask,
                                 o_icb_cmd_lock,
                                 o_icb_cmd_excl,
                                 o_icb_cmd_size_pre,
                                 o_icb_cmd_beat,
                                 o_icb_cmd_xlen_pre,
                                 o_icb_cmd_xburst,
                                 o_icb_cmd_modes,
                                 o_icb_cmd_dmode,
                                 o_icb_cmd_attri,
                                 o_icb_cmd_id,
                                 o_icb_cmd_usr} = cmd_fifo_o_dat;
  wire cmd_fifo_i_valid;
  wire cmd_fifo_i_ready;
  wire outs_cnt_full;
  assign cmd_fifo_i_valid = (~i_icb_reset_flag_r) & (~outs_cnt_full) & i_icb_cmd_valid;
  assign i_icb_cmd_ready  = (~i_icb_reset_flag_r) & (~outs_cnt_full) & cmd_fifo_i_ready;
  wire o_icb_cmd_valid_pre;
  wire o_icb_cmd_ready_pre;
  wire i_cmd_cdc_active;
  wire o_cmd_cdc_active;
  wire i_rsp_cdc_active;
  wire o_rsp_cdc_active;
  generate
  if(ASYNC_FIFO == 0) begin: cdc_buf_cmd
  e603_subsys_gnrl_cdc_buf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DW     (CMD_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_buf_cmd(
    .i_clk    (i_clk),
    .i_rst_n  (i_rst_n),
    .i_vld    (cmd_fifo_i_valid),
    .i_rdy    (cmd_fifo_i_ready),
    .i_dat    (cmd_fifo_i_dat),
    .i_cdc_buf_active(i_cmd_cdc_active),
    .o_cdc_buf_active(o_cmd_cdc_active),
    .o_clk    (o_clk),
    .o_rst_n  (o_rst_n),
    .o_vld    (o_icb_cmd_valid_pre),
    .o_rdy    (o_icb_cmd_ready_pre),
    .o_dat    (cmd_fifo_o_dat )
  );
  end
  else begin: cdc_fifo_cmd
  e603_subsys_gnrl_cdc_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (CMD_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_cmd(
    .i_clk    (i_clk),
    .i_rst_n  (i_rst_n),
    .i_vld    (cmd_fifo_i_valid),
    .i_rdy    (cmd_fifo_i_ready),
    .i_dat    (cmd_fifo_i_dat),
    .i_cdc_fifo_active(i_cmd_cdc_active),
    .o_cdc_fifo_active(o_cmd_cdc_active),
    .o_clk    (o_clk),
    .o_rst_n  (o_rst_n),
    .o_vld    (o_icb_cmd_valid_pre),
    .o_rdy    (o_icb_cmd_ready_pre),
    .o_dat    (cmd_fifo_o_dat )
  );
  end
  endgenerate
  wire o_outs_cnt_max;
  wire rsp_buf_ready;
  generate
    if(RSP_ALWAYS_READY == 1) begin: gen_rsp_always_ready_1
      assign o_icb_cmd_valid     = rsp_buf_ready & o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = rsp_buf_ready & o_icb_cmd_ready;
    end
    else begin: gen_rsp_always_ready_0
      assign o_icb_cmd_valid     = o_icb_cmd_valid_pre;
      assign o_icb_cmd_ready_pre = o_icb_cmd_ready;
    end
  endgenerate
  assign o_icb_cmd_sel = o_icb_cmd_valid_pre;
  localparam RSP_PACK_W = (2+DW+RSP_UW+ID_W+1+0);
  wire [RSP_PACK_W-1:0] rsp_fifo_i_dat = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata,
                                 o_icb_rsp_id,
                                 o_icb_rsp_last,
                                 o_icb_rsp_usr};
  wire [RSP_PACK_W-1:0] rsp_fifo_o_dat;
  assign {
                                 i_icb_rsp_err,
                                 i_icb_rsp_excl_ok,
                                 i_icb_rsp_rdata,
                                 i_icb_rsp_id,
                                 i_icb_rsp_last,
                                 i_icb_rsp_usr} = rsp_fifo_o_dat;
  wire o_icb_rsp_valid_raw;
  wire o_icb_rsp_ready_raw;
  generate
  if(ASYNC_FIFO == 0) begin: cdc_buf_rsp
  e603_subsys_gnrl_cdc_buf # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DW     (RSP_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_buf_rsp(
    .i_clk    (o_clk),
    .i_rst_n  (o_rst_n),
    .i_vld   (o_icb_rsp_valid_raw),
    .i_rdy   (o_icb_rsp_ready_raw),
    .i_dat   (rsp_fifo_i_dat ),
    .i_cdc_buf_active(o_rsp_cdc_active),
    .o_cdc_buf_active(i_rsp_cdc_active),
    .o_clk    (i_clk),
    .o_rst_n  (i_rst_n),
    .o_vld  (i_icb_rsp_valid),
    .o_rdy  (i_icb_rsp_ready),
    .o_dat  (rsp_fifo_o_dat )
  );
  end
  else begin: cdc_fifo_rsp
  e603_subsys_gnrl_cdc_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DP(ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (RSP_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_rsp(
    .i_clk    (o_clk),
    .i_rst_n  (o_rst_n),
    .i_vld   (o_icb_rsp_valid_raw),
    .i_rdy   (o_icb_rsp_ready_raw),
    .i_dat   (rsp_fifo_i_dat ),
    .i_cdc_fifo_active(o_rsp_cdc_active),
    .o_cdc_fifo_active(i_rsp_cdc_active),
    .o_clk    (i_clk),
    .o_rst_n  (i_rst_n),
    .o_vld  (i_icb_rsp_valid),
    .o_rdy  (i_icb_rsp_ready),
    .o_dat  (rsp_fifo_o_dat )
  );
  end
  endgenerate
  wire outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready
                    ;
  wire outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready
                    ;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] outs_cnt_r;
  wire [OUTS_CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, i_clk, i_rst_n);// VPP_NO_REG_PARSE
  assign outs_cnt_full = (outs_cnt_r == {OUTS_CNT_W{1'b1}});
  wire o_outs_cnt_inc = o_icb_cmd_valid & o_icb_cmd_ready 
                    ;
  wire o_outs_cnt_dec = o_icb_rsp_valid & o_icb_rsp_ready 
                    ;
  wire o_outs_cnt_ena = o_outs_cnt_inc ^ o_outs_cnt_dec;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_r;
  wire [OUTS_CNT_W-1:0] o_outs_cnt_nxt = o_outs_cnt_inc ? (o_outs_cnt_r + 1'b1) : (o_outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(OUTS_CNT_W) o_outs_cnt_dfflr (o_outs_cnt_ena, o_outs_cnt_nxt, o_outs_cnt_r, o_clk, o_rst_n);// VPP_NO_REG_PARSE
  assign icb2icb_async_i_active = i_cmd_cdc_active | i_rsp_cdc_active | i_icb_cmd_valid | (~(outs_cnt_r == {OUTS_CNT_W{1'b0}}));
  assign icb2icb_async_o_active = o_cmd_cdc_active | o_rsp_cdc_active | o_icb_cmd_valid_pre | (~(o_outs_cnt_r == {OUTS_CNT_W{1'b0}}));
  wire o_outs_cnt_eq0 = (o_outs_cnt_r == {OUTS_CNT_W{1'b0}});
  assign o_outs_cnt_max = (o_outs_cnt_r == {OUTS_CNT_W{1'b1}});
  generate
  if (RSP_STRICT_ORDER == 1) begin: rsp_strict_order_gen
      assign o_icb_rsp_valid_raw = (~o_outs_cnt_eq0) & o_icb_rsp_valid;
      assign o_icb_rsp_ready     = (~o_outs_cnt_eq0) & o_icb_rsp_ready_raw;
  end
  else begin: rsp_no_order_gen
      assign o_icb_rsp_valid_raw = o_icb_rsp_valid;
      assign o_icb_rsp_ready     = o_icb_rsp_ready_raw;
  end
  endgenerate
  assign rsp_buf_ready = (o_outs_cnt_r == {OUTS_CNT_W{1'b0}}) & o_icb_rsp_ready;
endmodule
module e603_subsys_gnrl_ficb_n2w_id # (
    parameter ID_W = 4,
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 64
) (
  input              i_icb_cmd_sel ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [ID_W-1:0] i_icb_cmd_id,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
    wire cmd_y_lo_hi;
    wire rsp_y_lo_hi;
    wire rsp_y_lo_hi_real;
    wire rsp_y_merged;
    wire i_icb_rsp_hasked = i_icb_rsp_valid & i_icb_rsp_ready;
    assign rsp_y_lo_hi_real = rsp_y_lo_hi;
    wire i_icb_cmd_hasked = i_icb_cmd_valid & i_icb_cmd_ready;
    wire n2w_fifo_wen = o_icb_cmd_valid & o_icb_cmd_ready;
    wire n2w_fifo_ren = o_icb_rsp_valid & o_icb_rsp_ready;
    wire n2w_fifo_i_ready;
    wire n2w_fifo_i_valid = n2w_fifo_wen;
    wire n2w_fifo_full    = (~n2w_fifo_i_ready);
    wire n2w_fifo_o_valid ;
    wire n2w_fifo_o_ready = n2w_fifo_ren;
    wire n2w_fifo_empty   = (~n2w_fifo_o_valid);
    wire cmd_y_merged;
  generate
  if (ZEROCYC_RSP == 1) begin:gen_0cyc_rsp_1
      e603_subsys_gnrl_bypbuf #(
              .PAYLOAD_NORST(PAYLOAD_NORST),
              .DP  (FIFO_OUTS_NUM),
              .DW  (2+ID_W
                   )
      )  u_n2w_bypbuf(
          .i_vld(n2w_fifo_i_valid),
          .i_rdy(n2w_fifo_i_ready),
          .i_dat({
              i_icb_cmd_id,cmd_y_lo_hi, cmd_y_merged
              } ),
          .o_dat({
              i_icb_rsp_id,rsp_y_lo_hi, rsp_y_merged
              } ),
          .o_vld(n2w_fifo_o_valid),
          .o_rdy(n2w_fifo_o_ready),
          .fifo_o_vld(),
          .clk(clk),
          .rst_n(rst_n)
      );
  end
  else begin :gen_0cyc_rsp_0
      e603_subsys_gnrl_fifo # (
              .PAYLOAD_NORST(PAYLOAD_NORST),
        .CUT_READY (FIFO_CUT_READY),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
              .DW  (2+ID_W
              )
      ) u_n2w_fifo (
        .i_vld(n2w_fifo_i_valid),
        .i_rdy(n2w_fifo_i_ready),
        .o_vld(n2w_fifo_o_valid),
        .o_rdy(n2w_fifo_o_ready),
          .i_dat({
              i_icb_cmd_id,cmd_y_lo_hi, cmd_y_merged
              } ),
          .o_dat({
              i_icb_rsp_id,rsp_y_lo_hi, rsp_y_merged
              } ),
        .clk  (clk),
        .rst_n(rst_n)
      );
  end
  endgenerate
  wire [AW-1:0]    i_icb_cmd_addr_algn;
  wire i_icb_cmd_size_full;
  wire i_icb_cmd_addr_lowr;
  generate
    if(X_W == 32) begin: gen_x_w_32
        assign cmd_y_lo_hi = i_icb_cmd_addr[2];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b10);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[2];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:3],3'b0};
    end
    if(X_W == 64) begin: gen_x_w_64
        assign cmd_y_lo_hi = i_icb_cmd_addr[3];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b11);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[3];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:4],4'b0};
    end
    if(X_W == 128) begin: gen_x_w_128
        assign cmd_y_lo_hi = i_icb_cmd_addr[4];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b100);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[4];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:5],5'b0};
    end
    if(X_W == 256) begin: gen_x_w_256
        assign cmd_y_lo_hi = i_icb_cmd_addr[5];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b101);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[5];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:6],6'b0};
    end
    if(X_W == 512) begin: gen_x_w_512
        assign cmd_y_lo_hi = i_icb_cmd_addr[6];
        assign i_icb_cmd_size_full = (i_icb_cmd_size[2:0] == 3'b110);
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[6];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:7],7'b0};
    end
    if(X_W == 1024) begin: gen_x_w_1024
        assign cmd_y_lo_hi = i_icb_cmd_addr[7];
        assign i_icb_cmd_size_full = 1'b0;
        assign i_icb_cmd_addr_lowr = ~i_icb_cmd_addr[7];
        assign i_icb_cmd_addr_algn = {i_icb_cmd_addr[AW-1:8],8'b0};
    end
  endgenerate
  wire icb_2nd_flag_r;
  wire i_icb_cmd_fixed = (i_icb_cmd_xburst == 2'b00);
  wire i_icb_cmd_wrap = (i_icb_cmd_xburst == 2'b10);
  wire i_icb_cmd_wrap_xlen1 = i_icb_cmd_wrap & (~(| i_icb_cmd_xlen[7:1])) & i_icb_cmd_xlen[0];
  wire   i_icb_cmd_need_merg_pre =                    
                       (i_icb_cmd_xlen[0]) & 
                       i_icb_cmd_size_full &
                       ( i_icb_cmd_wrap_xlen1 ? 1'b1 : 
                                                i_icb_cmd_addr_lowr 
                       )
                       & (~i_icb_cmd_fixed)
                       ;
  wire   i_icb_cmd_need_merg = (~icb_2nd_flag_r) & i_icb_cmd_need_merg_pre;
  wire [Y_W-1:0]     o_icb_cmd_wdata_pre;
  wire [(Y_W/8-1):0] o_icb_cmd_wmask_pre;
  assign o_icb_cmd_wdata_pre = {i_icb_cmd_wdata,i_icb_cmd_wdata};
  assign o_icb_cmd_wmask_pre = cmd_y_lo_hi ?  {i_icb_cmd_wmask,  {X_W/8{1'b0}}} : {  {X_W/8{1'b0}},i_icb_cmd_wmask};
  wire i_icb_cmd_xlen_is1 = (i_icb_cmd_xlen == 8'd1);
  wire i_icb_cmd_xlen_is0 = (i_icb_cmd_xlen == 8'd0);
  wire i_cmd_xlen_cvt_incr = i_icb_cmd_xlen_is1 & i_icb_cmd_need_merg_pre;
  wire icb_2nd_cmd_valid_r;
  wire icb_2nd_cmd_read_r;
  wire i_icb_cmd_read_need_merg = 1'b0;
  assign cmd_y_merged = ( icb_2nd_cmd_valid_r 
                        )
                        ;
  wire o_icb_cmd_hasked  = o_icb_cmd_valid & o_icb_cmd_ready;
  wire n2w_icb_2nd_cmd_valid_set_raw = i_icb_cmd_need_merg & (~icb_2nd_cmd_valid_r); 
  wire n2w_icb_2nd_cmd_valid_set = n2w_icb_2nd_cmd_valid_set_raw & i_icb_cmd_hasked
             ;
  wire icb_2nd_cmd_valid_clr = o_icb_cmd_hasked & icb_2nd_cmd_valid_r;
  wire icb_2nd_cmd_valid_ena = n2w_icb_2nd_cmd_valid_set | icb_2nd_cmd_valid_clr;
  wire icb_2nd_cmd_valid_nxt = n2w_icb_2nd_cmd_valid_set;
e603_subsys_gnrl_dfflr #(1) icb_2nd_cmd_valid (icb_2nd_cmd_valid_ena, icb_2nd_cmd_valid_nxt, icb_2nd_cmd_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_2nd_flag_set = (~i_icb_cmd_xlen_is0) & i_icb_cmd_hasked & (~icb_2nd_flag_r) & (~i_icb_cmd_beat[1]);
  wire icb_2nd_flag_clr = i_icb_cmd_hasked & icb_2nd_flag_r;
  wire icb_2nd_flag_ena = icb_2nd_flag_set | icb_2nd_flag_clr;
  wire icb_2nd_flag_nxt = (~icb_2nd_flag_clr);
e603_subsys_gnrl_dfflr #(1) icb_2nd_flag (icb_2nd_flag_ena, icb_2nd_flag_nxt, icb_2nd_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire merg_buf_ena = n2w_icb_2nd_cmd_valid_set;
  wire [AW-1:0]    icb_2nd_cmd_addr_r;
  wire [X_W-1:0]   icb_2nd_cmd_wdata_r;
  wire [X_W/8-1:0] icb_2nd_cmd_wmask_r;
  wire             icb_2nd_cmd_beat0_r;
  wire i_icb_cmd_beat0 = i_icb_cmd_beat[0] & (~i_icb_cmd_xlen_is1);
e603_subsys_gnrl_dffl  #(AW)   icb_2nd_cmd_addr (merg_buf_ena, i_icb_cmd_addr_algn , icb_2nd_cmd_addr_r , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(X_W)  icb_2nd_cmd_wdata(merg_buf_ena, i_icb_cmd_wdata, icb_2nd_cmd_wdata_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(X_W/8)icb_2nd_cmd_wmask(merg_buf_ena, i_icb_cmd_wmask, icb_2nd_cmd_wmask_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)    icb_2nd_cmd_beat0(merg_buf_ena, i_icb_cmd_beat0 , icb_2nd_cmd_beat0_r , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)    icb_2nd_cmd_read (merg_buf_ena, i_icb_cmd_read  , icb_2nd_cmd_read_r  , clk, rst_n);// VPP_NO_REG_PARSE
  assign o_icb_cmd_sel   = (~n2w_fifo_full) & (i_icb_cmd_sel   | icb_2nd_cmd_valid_r);
  assign o_icb_cmd_valid = (~n2w_fifo_full) & (i_icb_cmd_need_merg ? (i_icb_cmd_valid & icb_2nd_cmd_valid_r) : i_icb_cmd_valid);
  assign i_icb_cmd_ready = (~n2w_fifo_full) & ((i_icb_cmd_need_merg & (~icb_2nd_cmd_valid_r)) ? 1'b1 : o_icb_cmd_ready);
  assign o_icb_cmd_addr  = 
            icb_2nd_cmd_valid_r ? icb_2nd_cmd_addr_r : i_icb_cmd_addr;
  assign o_icb_cmd_wdata = icb_2nd_cmd_valid_r ? (
                                 cmd_y_lo_hi ? {i_icb_cmd_wdata, icb_2nd_cmd_wdata_r} : {icb_2nd_cmd_wdata_r, i_icb_cmd_wdata}
                                 ) : o_icb_cmd_wdata_pre;
  assign o_icb_cmd_wmask = icb_2nd_cmd_valid_r ? (
                                 cmd_y_lo_hi ? {i_icb_cmd_wmask, icb_2nd_cmd_wmask_r} : {icb_2nd_cmd_wmask_r, i_icb_cmd_wmask}
                                 ) : o_icb_cmd_wmask_pre;
  wire             o_icb_cmd_read_pre;
  wire             o_icb_cmd_lock_pre;
  wire             o_icb_cmd_excl_pre;
  wire [1:0]       o_icb_cmd_modes_pre;
  wire             o_icb_cmd_dmode_pre;
  wire [1:0]       o_icb_cmd_xburst_pre;
  wire [2:0]       o_icb_cmd_attri_pre;
  assign o_icb_cmd_read_pre   = i_icb_cmd_read;
  assign o_icb_cmd_lock_pre   = i_icb_cmd_lock;
  assign o_icb_cmd_excl_pre   = i_icb_cmd_excl;
  assign o_icb_cmd_usr    = i_icb_cmd_usr;
  wire [ID_W-1:0] o_icb_cmd_id_pre;
  assign o_icb_cmd_id_pre    = {ID_W{1'b0}};
  assign o_icb_cmd_id = o_icb_cmd_id_pre;
  assign o_icb_cmd_xburst_pre = i_cmd_xlen_cvt_incr ? 2'b01 : i_icb_cmd_xburst;
  assign o_icb_cmd_modes_pre  = i_icb_cmd_modes ;
  assign o_icb_cmd_dmode_pre  = i_icb_cmd_dmode ;
  assign o_icb_cmd_attri_pre  = i_icb_cmd_attri ;
  assign o_icb_cmd_read   = o_icb_cmd_read_pre;
  assign o_icb_cmd_lock   = o_icb_cmd_lock_pre;
  assign o_icb_cmd_excl   = o_icb_cmd_excl_pre;
  assign o_icb_cmd_modes  = o_icb_cmd_modes_pre;
  assign o_icb_cmd_dmode  = o_icb_cmd_dmode_pre;
  assign o_icb_cmd_xburst = o_icb_cmd_xburst_pre;
  assign o_icb_cmd_attri  = o_icb_cmd_attri_pre;
  wire [2:0] o_icb_cmd_size_pre;
  wire [7:0] o_icb_cmd_xlen_pre;
  wire [1:0] o_icb_cmd_beat_pre;
  assign o_icb_cmd_size = o_icb_cmd_size_pre;
  assign o_icb_cmd_xlen = o_icb_cmd_xlen_pre;
  assign o_icb_cmd_beat = o_icb_cmd_beat_pre;
  assign o_icb_cmd_beat_pre[0] = (icb_2nd_cmd_valid_r ? icb_2nd_cmd_beat0_r : i_icb_cmd_beat[0]) & (~i_cmd_xlen_cvt_incr);
  assign o_icb_cmd_beat_pre[1] = i_icb_cmd_beat[1] & (~(icb_2nd_cmd_valid_r & i_icb_cmd_xlen_is1));
  generate
  if (X_W == 32) begin:dw_64_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b011 : i_icb_cmd_size;
  end
  if (X_W == 64) begin:dw_128_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b100 : i_icb_cmd_size;
  end
  if (X_W == 128) begin:dw_256_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b101 : i_icb_cmd_size;
  end
  if (X_W == 256) begin:dw_512_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b110 : i_icb_cmd_size;
  end
  if (X_W == 512) begin:dw_1024_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b111 : i_icb_cmd_size;
  end
  if (X_W == 1024) begin:dw_2048_o_icb
    assign o_icb_cmd_size_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? 3'b111 : i_icb_cmd_size;
  end
  endgenerate
    assign o_icb_cmd_xlen_pre = (icb_2nd_cmd_valid_r | i_icb_cmd_read_need_merg) ? {1'b0,i_icb_cmd_xlen[7:1]} : i_icb_cmd_xlen;
  wire icb_2nd_rsp_valid_r;
  wire icb_2nd_rsp_valid_set = (~icb_2nd_rsp_valid_r) & rsp_y_merged & i_icb_rsp_hasked;
  wire icb_2nd_rsp_valid_clr = icb_2nd_rsp_valid_r & i_icb_rsp_hasked;
  wire icb_2nd_rsp_valid_ena = icb_2nd_rsp_valid_set | icb_2nd_rsp_valid_clr;
  wire icb_2nd_rsp_valid_nxt = icb_2nd_rsp_valid_set;
e603_subsys_gnrl_dfflr #(1) icb_2nd_rsp_valid (icb_2nd_rsp_valid_ena, icb_2nd_rsp_valid_nxt, icb_2nd_rsp_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign o_icb_rsp_ready = (rsp_y_merged ? icb_2nd_rsp_valid_r : 1'b1) & i_icb_rsp_ready & n2w_fifo_o_valid;
  wire [X_W-1:0] i_icb_rsp_rdata_pre;
  wire [X_W-1:0] i_icb_rsp_rdata_merged;
  assign i_icb_rsp_rdata_pre    = rsp_y_lo_hi_real ? o_icb_rsp_rdata[Y_W-1:X_W] : o_icb_rsp_rdata[X_W-1:0] ;
  wire i_icb_rsp_rdata_merged_sel = (icb_2nd_rsp_valid_r ? rsp_y_lo_hi : (~rsp_y_lo_hi)); 
  assign i_icb_rsp_rdata_merged = i_icb_rsp_rdata_merged_sel 
                                     ? o_icb_rsp_rdata[Y_W-1:X_W] : o_icb_rsp_rdata[X_W-1:0] ;
  assign i_icb_rsp_rdata = rsp_y_merged ? i_icb_rsp_rdata_merged : i_icb_rsp_rdata_pre;
  assign i_icb_rsp_valid   = o_icb_rsp_valid & n2w_fifo_o_valid;  
  assign i_icb_rsp_err     = o_icb_rsp_err   ;
  assign i_icb_rsp_excl_ok = o_icb_rsp_excl_ok   ;
  assign i_icb_rsp_usr   = o_icb_rsp_usr   ;
  assign i_icb_rsp_last   = rsp_y_merged ? (icb_2nd_rsp_valid_r & o_icb_rsp_last)  :  o_icb_rsp_last;
endmodule
module e603_subsys_gnrl_ficb_nn2ww_id # (
    parameter ID_W = 4,
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 128
) (
  input              i_icb_cmd_sel ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [ID_W-1:0] i_icb_cmd_id,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel  ,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W*2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W/4-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [ID_W-1:0]  dw_icb_cmd_id;
  wire [7:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W*2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
  wire [ID_W-1:0]  dw_icb_rsp_id;
  wire             dw_icb_rsp_last;
  e603_subsys_gnrl_ficb_n2w_id # (
    .ID_W(ID_W),
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W*2 )
  ) u_ficb_32to64 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id       (i_icb_cmd_id    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id       (i_icb_rsp_id    ),
    .i_icb_rsp_last       (i_icb_rsp_last    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel   ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_id       (dw_icb_cmd_id     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .o_icb_rsp_id       (dw_icb_rsp_id     ),
    .o_icb_rsp_last       (dw_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_n2w_id # (
    .ID_W(ID_W),
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W*2),
    .Y_W(Y_W )
  ) u_ficb_64to128 (
    .i_icb_cmd_sel       (dw_icb_cmd_sel  ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_id       (dw_icb_cmd_id    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .i_icb_rsp_id       (dw_icb_rsp_id    ),
    .i_icb_rsp_last       (dw_icb_rsp_last    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id       (o_icb_cmd_id     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id       (o_icb_rsp_id     ),
    .o_icb_rsp_last       (o_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_nnn2www_id # (
    parameter ID_W = 4,
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 32,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 128
) (
  input              i_icb_cmd_sel ,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [ID_W-1:0] i_icb_cmd_id,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel  ,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W*2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W*2/8-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [ID_W-1:0]  dw_icb_cmd_id;
  wire [7:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W*2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
  wire [ID_W-1:0]  dw_icb_rsp_id;
  wire             dw_icb_rsp_last;
  wire               dw2_icb_cmd_sel;
  wire               dw2_icb_cmd_valid;
  wire               dw2_icb_cmd_ready;
  wire               dw2_icb_cmd_read;
  wire [AW-1:0]      dw2_icb_cmd_addr;
  wire [X_W*4-1:0]      dw2_icb_cmd_wdata;
  wire [(X_W*4/8-1):0]  dw2_icb_cmd_wmask;
  wire               dw2_icb_cmd_lock;
  wire               dw2_icb_cmd_excl;
  wire [2:0]         dw2_icb_cmd_size;
  wire [1:0]         dw2_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw2_icb_cmd_usr;
  wire [ID_W-1:0]  dw2_icb_cmd_id;
  wire [7:0]         dw2_icb_cmd_xlen;
  wire [1:0]         dw2_icb_cmd_xburst;
  wire [1:0]         dw2_icb_cmd_modes;
  wire               dw2_icb_cmd_dmode;
  wire [2:0]         dw2_icb_cmd_attri;
  wire               dw2_icb_rsp_valid;
  wire               dw2_icb_rsp_ready;
  wire               dw2_icb_rsp_err;
  wire               dw2_icb_rsp_excl_ok;
  wire [X_W*4-1:0]      dw2_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw2_icb_rsp_usr;
  wire [ID_W-1:0]  dw2_icb_rsp_id;
  wire             dw2_icb_rsp_last;
  e603_subsys_gnrl_ficb_n2w_id # (
    .ID_W(ID_W),
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W*2 )
  ) u_ficb_x_to_xm2 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id       (i_icb_cmd_id    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id       (i_icb_rsp_id    ),
    .i_icb_rsp_last       (i_icb_rsp_last    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel   ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_id       (dw_icb_cmd_id     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .o_icb_rsp_id       (dw_icb_rsp_id     ),
    .o_icb_rsp_last       (dw_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_n2w_id # (
    .ID_W(ID_W),
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W*2),
    .Y_W(X_W*4)
  ) u_ficb_xm2_to_xm4 (
    .i_icb_cmd_sel       (dw_icb_cmd_sel  ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_id       (dw_icb_cmd_id    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .i_icb_rsp_id       (dw_icb_rsp_id    ),
    .i_icb_rsp_last       (dw_icb_rsp_last    ),
    .o_icb_cmd_sel       (dw2_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw2_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw2_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw2_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw2_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw2_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw2_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw2_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw2_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw2_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw2_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw2_icb_cmd_usr     ),
    .o_icb_cmd_id       (dw2_icb_cmd_id     ),
    .o_icb_cmd_xlen      (dw2_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw2_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw2_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw2_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw2_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw2_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw2_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw2_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw2_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw2_icb_rsp_usr     ),
    .o_icb_rsp_id       (dw2_icb_rsp_id     ),
    .o_icb_rsp_last       (dw2_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_n2w_id # (
    .ID_W(ID_W),
    .PAYLOAD_NORST   (PAYLOAD_NORST   ),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W*4),
    .Y_W(Y_W)
  ) u_ficb_xm4_to_y (
    .i_icb_cmd_sel       (dw2_icb_cmd_sel  ),
    .i_icb_cmd_valid     (dw2_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw2_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw2_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw2_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw2_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw2_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw2_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw2_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw2_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw2_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw2_icb_cmd_usr    ),
    .i_icb_cmd_id       (dw2_icb_cmd_id    ),
    .i_icb_cmd_xlen      (dw2_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw2_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw2_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw2_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw2_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw2_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw2_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw2_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw2_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw2_icb_rsp_usr    ),
    .i_icb_rsp_id       (dw2_icb_rsp_id    ),
    .i_icb_rsp_last       (dw2_icb_rsp_last    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id       (o_icb_cmd_id     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id       (o_icb_rsp_id     ),
    .o_icb_rsp_last       (o_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_w2n_id # (
    parameter ID_W = 4,
    parameter FIFO_OUTS_CNT_W = 3,
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 1,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 64,
  parameter Y_W = 32
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [ID_W-1:0] i_icb_cmd_id,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  wire i_icb_rsp_err_pre;
  wire i_icb_rsp_excl_ok_pre;
  assign i_icb_rsp_err = i_icb_rsp_err_pre;
  assign i_icb_rsp_excl_ok = i_icb_rsp_excl_ok_pre;
  wire icb_cmd_size_dw;
  wire icb_cmd_addr_2 ;
  wire icb_cmd_size_dw_real = icb_cmd_size_dw;
generate
if (X_W == 64) begin:dw_64
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b11);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[2];
end
if (X_W == 128) begin:dw_128
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b100);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[3];
end
if (X_W == 256) begin:dw_256
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b101);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[4];
end
if (X_W == 512) begin:dw_512
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b110);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[5];
end
if (X_W == 1024) begin:dw_1024
  assign icb_cmd_size_dw = (i_icb_cmd_size[2:0] == 3'b111);
  assign icb_cmd_addr_2  = i_icb_cmd_addr[6];
end
endgenerate
  wire o_icb_rsp_hasked  = o_icb_rsp_valid & o_icb_rsp_ready;
    wire icb_rsp_fixed_cvt;
    wire icb_rsp_write;
wire i_icb_cmd_fixed_cvt;
  wire w2n_fifo_wen = i_icb_cmd_valid & i_icb_cmd_ready;
  wire w2n_fifo_ren = i_icb_rsp_valid & i_icb_rsp_ready;
  wire w2n_fifo_i_valid = w2n_fifo_wen;
  wire w2n_fifo_i_ready;
  wire w2n_fifo_o_valid;
  wire w2n_fifo_o_match;
  wire w2n_has_ooo_id_buf;
  wire w2n_fifo_o_ready = w2n_fifo_ren;
  wire w2n_fifo_full;
    wire i_icb_cmd_xlen_is0 = (i_icb_cmd_xlen == {O_AXLEN_W{1'b0}});
    wire i_icb_xlen_overflow;
    wire icb_2nd_xlen_overflow;
    wire i_icb_cmd_xburst_fixed = (i_icb_cmd_xburst[1:0] == 2'b0);
    wire i_icb_cmd_xburst_fixed_xlen0     = (i_icb_cmd_xlen_is0 & i_icb_cmd_xburst_fixed);
    wire i_icb_cmd_xburst_fixed_n_xlen0 = ((~i_icb_cmd_xlen_is0) & i_icb_cmd_xburst_fixed);
    wire [1:0] i_icb_cmd_xburst_cvt = (i_icb_cmd_xburst_fixed_xlen0) ? 2'b01 : i_icb_cmd_xburst[1:0];
    assign i_icb_cmd_fixed_cvt = i_icb_cmd_xburst_fixed_n_xlen0 | i_icb_xlen_overflow; 
  wire icb_rsp_size_dw;
  wire icb_2nd_rsp_valid_r;
  wire o_icb_rsp_valid_dw = (icb_rsp_size_dw ? icb_2nd_rsp_valid_r : 1'b1);
generate
if(SUPPORT_W2N_ID_OOO == 1) begin: id_ooo_is1_full
  wire fixed_outs_cnt_inc = i_icb_cmd_valid & i_icb_cmd_ready & i_icb_cmd_fixed_cvt;
  wire fixed_outs_cnt_dec = i_icb_rsp_valid & i_icb_rsp_ready & icb_rsp_fixed_cvt;
  wire fixed_outs_cnt_ena = fixed_outs_cnt_inc ^ fixed_outs_cnt_dec;
  wire [FIFO_OUTS_CNT_W-1:0] fixed_outs_cnt_r;
  wire [FIFO_OUTS_CNT_W-1:0] fixed_outs_cnt_nxt = fixed_outs_cnt_inc ? (fixed_outs_cnt_r + 1'b1) : (fixed_outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(FIFO_OUTS_CNT_W)         fixed_outs_cnt_dfflr (fixed_outs_cnt_ena, fixed_outs_cnt_nxt, fixed_outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire fixed_outs_cnt_eq0 = (fixed_outs_cnt_r == {{FIFO_OUTS_CNT_W-1{1'b0}},1'b0});
  wire any_fixed_outstanding = ~fixed_outs_cnt_eq0; 
  assign w2n_fifo_full = (~w2n_fifo_i_ready) | any_fixed_outstanding 
                       | (w2n_fifo_o_valid & i_icb_cmd_fixed_cvt);
end
else begin: id_ooo_is0_full
  assign w2n_fifo_full = ~w2n_fifo_i_ready;
end
endgenerate
  wire w2n_fifo_empty = ~w2n_fifo_o_valid;
  wire icb_rsp_addr_2;
  wire icb_2nd_cmd_read_r;
  wire i_icb_cmd_last = i_icb_cmd_beat[1] | (i_icb_cmd_xlen == {O_AXLEN_W{1'b0}});
    wire icb_cmd_last = i_icb_cmd_last;
    wire icb_rsp_last;
generate
if (ZEROCYC_RSP == 1) begin:gen_0cyc_rsp_1
    assign w2n_has_ooo_id_buf = 1'b0;
    assign w2n_fifo_o_match = 1'b0;
  e603_subsys_gnrl_bypbuf #(
    .PAYLOAD_NORST(PAYLOAD_NORST),
          .DP  (FIFO_OUTS_NUM),
          .DW  (2+ID_W+1
               )
  )  u_rsp_w2n_bypbuf(
      .i_vld(w2n_fifo_i_valid),
      .i_rdy(w2n_fifo_i_ready),
      .i_dat({
              i_icb_cmd_id, i_icb_cmd_last, icb_cmd_size_dw_real,icb_cmd_addr_2
              }),
      .o_dat({
              i_icb_rsp_id, i_icb_rsp_last, icb_rsp_size_dw,icb_rsp_addr_2
              }),
      .o_vld(w2n_fifo_o_valid),
      .o_rdy(w2n_fifo_o_ready),
      .fifo_o_vld(),
      .clk(clk),
      .rst_n(rst_n)
  );
end
else begin :gen_0cyc_rsp_0
    if(SUPPORT_W2N_ID_OOO == 1) begin: id_ooo_is1
    assign w2n_has_ooo_id_buf = 1'b1;
      e603_subsys_ficbw2n_gnrl_ooo_id_buf # (
        .IDW(ID_W),
        .DP_PTR_W(FIFO_OUTS_CNT_W),
          .DW  (4
          ),
          .DP  (FIFO_OUTS_NUM) 
      )  u_rsp_w2n_fifo(
          .i_vld(w2n_fifo_i_valid),
          .i_rdy(w2n_fifo_i_ready),
          .i_dat({i_icb_cmd_fixed_cvt,icb_cmd_last,icb_cmd_size_dw_real,icb_cmd_addr_2
          }),
          .o_dat({icb_rsp_fixed_cvt,icb_rsp_last,icb_rsp_size_dw,icb_rsp_addr_2
          }),
        .i_id(i_icb_cmd_id),
        .o_id(i_icb_rsp_id),
          .o_match(w2n_fifo_o_match),
          .o_vld(w2n_fifo_o_valid),
          .o_rdy(w2n_fifo_o_ready),
          .clk(clk),
          .rst_n(rst_n)
      );
    end
    else begin: id_ooo_is0
    assign w2n_has_ooo_id_buf = 1'b0;
    assign w2n_fifo_o_match = 1'b0;
      e603_subsys_gnrl_fifo #(
    .PAYLOAD_NORST(PAYLOAD_NORST),
          .CUT_READY (FIFO_CUT_READY),
          .MSKO      (0),
          .DP  (FIFO_OUTS_NUM),
          .DW  (2+ID_W+1 
             )
      )  u_rsp_w2n_fifo(
          .i_vld(w2n_fifo_i_valid),
          .i_rdy(w2n_fifo_i_ready),
      .i_dat({
              i_icb_cmd_id, i_icb_cmd_last, icb_cmd_size_dw_real,icb_cmd_addr_2
              }),
      .o_dat({
              i_icb_rsp_id, i_icb_rsp_last, icb_rsp_size_dw,icb_rsp_addr_2
              }),
          .o_vld(w2n_fifo_o_valid),
          .o_rdy(w2n_fifo_o_ready),
          .clk(clk),
          .rst_n(rst_n)
      );
    end
end
endgenerate
  wire             icb_2nd_cmd_valid_r;
  wire             icb_2nd_cmd_valid_ena;
  wire             icb_2nd_cmd_valid_nxt;
  wire             icb_2nd_cmd_valid_set;
  wire             icb_2nd_cmd_valid_clr;
  wire             i_icb_cmd_ready_addi_cond;
  wire o_icb_cmd_hasked  = o_icb_cmd_valid & o_icb_cmd_ready;
    wire i_icb_cvt_single;
    wire icb_2nd_cmd_valid_set_raw     = icb_cmd_size_dw      & o_icb_cmd_hasked & (~icb_2nd_cmd_valid_r);
    assign icb_2nd_cmd_valid_set     = icb_2nd_cmd_valid_set_raw;
    wire icb_2nd_cmd_set = icb_2nd_cmd_valid_set;
    assign icb_2nd_cmd_valid_clr     = icb_2nd_cmd_valid_r  & o_icb_cmd_hasked;
    wire icb_2nd_cmd_valid_real;
    assign icb_2nd_cmd_valid_real = icb_2nd_cmd_valid_r;
    assign i_icb_cmd_ready_addi_cond = !icb_2nd_cmd_valid_real;
    assign i_icb_cmd_ready = (~w2n_fifo_full) & i_icb_cmd_ready_addi_cond & o_icb_cmd_ready;
    wire             icb_2nd_cmd_excl_r;
    wire             icb_2nd_cmd_lock_r;
    wire [AW-1:0]    icb_2nd_cmd_addr_r;
    wire [Y_W-1:0]   icb_2nd_cmd_wdata_r;
    wire [Y_W/8-1:0] icb_2nd_cmd_wmask_r;
    wire [CMD_UW-1:0] icb_2nd_cmd_usr_r;
    wire [ID_W-1:0] icb_2nd_cmd_id_r;
    wire [1:0] icb_2nd_cmd_beat_r;
    wire [O_AXLEN_W-1:0] icb_2nd_cmd_xlen_r  ;
    wire [1:0] icb_2nd_cmd_xburst_r;
    wire [1:0] icb_2nd_cmd_modes_r ;
    wire icb_2nd_load_ena = icb_2nd_cmd_set;
    wire       icb_2nd_cmd_dmode_r ;
    wire [2:0] icb_2nd_cmd_attri_r ;
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_lock   (icb_2nd_load_ena, i_icb_cmd_lock, icb_2nd_cmd_lock_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_excl   (icb_2nd_load_ena, i_icb_cmd_excl, icb_2nd_cmd_excl_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_read   (icb_2nd_load_ena, i_icb_cmd_read, icb_2nd_cmd_read_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(AW)  icb_2nd_cmd_addr   (icb_2nd_cmd_set, i_icb_cmd_addr[AW-1:0], icb_2nd_cmd_addr_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(Y_W)   icb_2nd_cmd_wdata  (icb_2nd_load_ena, i_icb_cmd_wdata[X_W-1:Y_W], icb_2nd_cmd_wdata_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(Y_W/8) icb_2nd_cmd_wmask  (icb_2nd_load_ena, i_icb_cmd_wmask[X_W/8-1:Y_W/8], icb_2nd_cmd_wmask_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(CMD_UW)icb_2nd_cmd_usr    (icb_2nd_load_ena, i_icb_cmd_usr, icb_2nd_cmd_usr_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(ID_W)icb_2nd_cmd_id    (icb_2nd_load_ena, i_icb_cmd_id, icb_2nd_cmd_id_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2)     icb_2nd_cmd_beat   (icb_2nd_load_ena, i_icb_cmd_beat, icb_2nd_cmd_beat_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(O_AXLEN_W)     icb_2nd_cmd_xlen   (icb_2nd_load_ena, i_icb_cmd_xlen  , icb_2nd_cmd_xlen_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2)     icb_2nd_cmd_xburst (icb_2nd_load_ena, i_icb_cmd_xburst_cvt, icb_2nd_cmd_xburst_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2)     icb_2nd_cmd_modes  (icb_2nd_load_ena, i_icb_cmd_modes , icb_2nd_cmd_modes_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(1)     icb_2nd_cmd_dmode  (icb_2nd_load_ena, i_icb_cmd_dmode , icb_2nd_cmd_dmode_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(3)     icb_2nd_cmd_attri  (icb_2nd_load_ena, i_icb_cmd_attri , icb_2nd_cmd_attri_r, clk, rst_n);// VPP_NO_REG_PARSE
    assign o_icb_cmd_sel   = (~w2n_fifo_full) & i_icb_cmd_sel   || icb_2nd_cmd_valid_real;
    assign o_icb_cmd_valid = (~w2n_fifo_full) & i_icb_cmd_valid || icb_2nd_cmd_valid_real;
  wire [2:0] o_icb_cmd_size_pre;
  wire [O_AXLEN_W-1:0] o_icb_cmd_xlen_pre;
  wire [1:0] o_icb_cmd_beat_pre;
  wire [AW-1:0] o_icb_cmd_addr_pre;
  assign o_icb_cmd_size = o_icb_cmd_size_pre;
  assign o_icb_cmd_xlen = o_icb_cmd_xlen_pre;
  assign o_icb_cmd_beat = o_icb_cmd_beat_pre;
  assign o_icb_cmd_addr = o_icb_cmd_addr_pre;
  wire             o_icb_cmd_read_pre;
  wire             o_icb_cmd_lock_pre;
  wire             o_icb_cmd_excl_pre;
  wire [1:0]       o_icb_cmd_modes_pre;
  wire             o_icb_cmd_dmode_pre;
  wire [1:0]       o_icb_cmd_xburst_pre;
  wire [2:0]       o_icb_cmd_attri_pre;
  assign o_icb_cmd_read   = o_icb_cmd_read_pre;
  assign o_icb_cmd_lock   = o_icb_cmd_lock_pre;
  assign o_icb_cmd_excl   = o_icb_cmd_excl_pre;
  assign o_icb_cmd_modes  = o_icb_cmd_modes_pre ;
  assign o_icb_cmd_dmode  = o_icb_cmd_dmode_pre ;
  assign o_icb_cmd_attri  = o_icb_cmd_attri_pre ;
  assign o_icb_cmd_xburst = o_icb_cmd_xburst_pre ;
    assign o_icb_cmd_addr_pre = icb_2nd_cmd_valid_r ? (
                                                    (X_W == 64) ? {icb_2nd_cmd_addr_r[AW-1:3],3'b100} :
                                                    (X_W == 256) ? {icb_2nd_cmd_addr_r[AW-1:5],5'b10000} :
                                                    (X_W == 512) ? {icb_2nd_cmd_addr_r[AW-1:6],6'b100000} :
                                                    (X_W == 1024) ? {icb_2nd_cmd_addr_r[AW-1:7],7'b1000000} :
                                                                  {icb_2nd_cmd_addr_r[AW-1:4],4'b1000}
                                                    ) :
                             icb_cmd_size_dw    ? (
                                                    (X_W == 64) ? {i_icb_cmd_addr[AW-1:3],3'b0} :
                                                    (X_W == 256) ? {i_icb_cmd_addr[AW-1:5],5'b0} :
                                                    (X_W == 512) ? {i_icb_cmd_addr[AW-1:6],6'b0} :
                                                    (X_W == 1024) ? {i_icb_cmd_addr[AW-1:7],7'b0} :
                                                                  {i_icb_cmd_addr[AW-1:4],4'b0}
                                                    )
                                                :  i_icb_cmd_addr;
    assign o_icb_cmd_read_pre = icb_2nd_cmd_valid_real ? icb_2nd_cmd_read_r
                                                : i_icb_cmd_read;
    assign o_icb_cmd_lock_pre = icb_2nd_cmd_valid_real ? icb_2nd_cmd_lock_r
                                                : i_icb_cmd_lock;
    assign o_icb_cmd_excl_pre = icb_2nd_cmd_valid_real ? icb_2nd_cmd_excl_r
                                                : i_icb_cmd_excl;
    assign o_icb_cmd_wdata = icb_2nd_cmd_valid_real ? icb_2nd_cmd_wdata_r :
                             icb_cmd_size_dw     ? i_icb_cmd_wdata[Y_W-1:0] :
                             icb_cmd_addr_2      ? i_icb_cmd_wdata[X_W-1:Y_W] :
                                                   i_icb_cmd_wdata[Y_W-1:0];
    assign o_icb_cmd_wmask = icb_2nd_cmd_valid_real ? icb_2nd_cmd_wmask_r :
                             icb_cmd_size_dw     ? i_icb_cmd_wmask[(Y_W/8-1):0] :
                             icb_cmd_addr_2      ? i_icb_cmd_wmask[(X_W/8-1):(Y_W/8)] :
                                                   i_icb_cmd_wmask[(Y_W/8-1):0];
    assign o_icb_cmd_usr  = icb_2nd_cmd_valid_real ? icb_2nd_cmd_usr_r : i_icb_cmd_usr;
  generate
    if(SUPPORT_W2N_ID_OOO == 1) begin: cmd_id_ooo_is1
        assign o_icb_cmd_id  = icb_2nd_cmd_valid_real ? icb_2nd_cmd_id_r : i_icb_cmd_id;
    end
    else begin: cmd_id_ooo_is0
        assign o_icb_cmd_id  = {ID_W{1'b0}};
    end
  endgenerate
  generate
    if(O_AXLEN_EXTEND == 1) begin: xlen_extend_1_gen
        assign i_icb_xlen_overflow   = 1'b0;
        assign icb_2nd_xlen_overflow = 1'b0;
    end
    else begin: xlen_extend_0_gen
        assign i_icb_xlen_overflow = 
                    (icb_cmd_size_dw & (i_icb_cmd_xburst == 2'b10)) ? i_icb_cmd_xlen[3] : 
                    (icb_cmd_size_dw & (i_icb_cmd_xburst == 2'b01)) ? i_icb_cmd_xlen[7] : 1'b0 ;
        assign icb_2nd_xlen_overflow= (
                   (icb_2nd_cmd_xburst_r == 2'b10) ? icb_2nd_cmd_xlen_r[3] :
                   (icb_2nd_cmd_xburst_r == 2'b01) ? icb_2nd_cmd_xlen_r[7] : 1'b0) ;
    end
  endgenerate
    wire icb_2nd_cvt_single = (icb_2nd_cmd_xburst_r == 2'b0) | icb_2nd_xlen_overflow;
    assign i_icb_cvt_single   = i_icb_cmd_fixed_cvt;
    wire icb_2nd_cmd_xlen_is0 = (icb_2nd_cmd_xlen_r == {O_AXLEN_W{1'd0}});
    assign o_icb_cmd_beat_pre[0] = icb_2nd_cmd_valid_r ? (1'b0                                                                    ) : ((~i_icb_cvt_single) & (i_icb_cmd_beat[0] | (icb_cmd_size_dw & i_icb_cmd_xlen_is0)));
    assign o_icb_cmd_beat_pre[1] = icb_2nd_cmd_valid_r ? ((~icb_2nd_cvt_single) & (icb_2nd_cmd_beat_r[1] | (icb_2nd_cmd_xlen_is0))) : ((~i_icb_cvt_single) & (icb_cmd_size_dw ? 1'b0 : i_icb_cmd_beat[1]));
    wire [O_AXLEN_W-1:0] o_icb_cmd_xlen_raw;
    generate
    if (X_W == 64) begin:dw_64_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b10 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 128) begin:dw_128_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b11 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 256) begin:dw_256_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b100: i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 512) begin:dw_512_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b101 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    if (X_W == 1024) begin:dw_1024_o_icb
      assign o_icb_cmd_size_pre = 
               (icb_cmd_size_dw || icb_2nd_cmd_valid_real)  ? 3'b110 : i_icb_cmd_size;
      assign o_icb_cmd_xlen_raw = icb_2nd_cmd_valid_real ? ({O_AXLEN_W{~icb_2nd_cvt_single}} & {icb_2nd_cmd_xlen_r[O_AXLEN_W-2:0],1'b1}) : ( {O_AXLEN_W{~i_icb_cvt_single}} & (icb_cmd_size_dw ? {i_icb_cmd_xlen[O_AXLEN_W-2:0],1'b1} : i_icb_cmd_xlen));
    end
    endgenerate
    assign o_icb_cmd_xlen_pre = o_icb_cmd_xlen_raw;
    assign o_icb_cmd_xburst_pre  = icb_2nd_cmd_valid_real ? (icb_2nd_cvt_single ? 2'b01 : icb_2nd_cmd_xburst_r)
                                                   : (i_icb_cvt_single ? 2'b01 : i_icb_cmd_xburst_cvt);
    assign o_icb_cmd_modes_pre   = icb_2nd_cmd_valid_real ? icb_2nd_cmd_modes_r  : i_icb_cmd_modes ;
    assign o_icb_cmd_dmode_pre   = icb_2nd_cmd_valid_real ? icb_2nd_cmd_dmode_r  : i_icb_cmd_dmode ;
    assign o_icb_cmd_attri_pre   = icb_2nd_cmd_valid_real ? icb_2nd_cmd_attri_r  : i_icb_cmd_attri ;
  assign icb_2nd_cmd_valid_ena = icb_2nd_cmd_valid_set | icb_2nd_cmd_valid_clr;
  assign icb_2nd_cmd_valid_nxt = icb_2nd_cmd_valid_set & (~icb_2nd_cmd_valid_clr);
e603_subsys_gnrl_dfflr #(1)     icb_2nd_cmd_valid  (icb_2nd_cmd_valid_ena, icb_2nd_cmd_valid_nxt, icb_2nd_cmd_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire i_icb_rsp_hasked  = i_icb_rsp_valid & i_icb_rsp_ready;
  wire icb_2nd_rsp_valid_set = icb_rsp_size_dw & o_icb_rsp_hasked & (~icb_2nd_rsp_valid_r);
  wire icb_2nd_rsp_valid_clr = icb_rsp_size_dw & o_icb_rsp_hasked & icb_2nd_rsp_valid_r;
  wire icb_2nd_rsp_valid_ena = icb_2nd_rsp_valid_set | icb_2nd_rsp_valid_clr;
  wire icb_2nd_rsp_valid_nxt = icb_2nd_rsp_valid_set & (~icb_2nd_rsp_valid_clr);
e603_subsys_gnrl_dfflr #(1) icb_2nd_rsp_valid_dfflr(icb_2nd_rsp_valid_ena, icb_2nd_rsp_valid_nxt, icb_2nd_rsp_valid_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_ena = icb_rsp_size_dw &  o_icb_rsp_hasked & (~icb_2nd_rsp_valid_r);
  wire [Y_W-1:0] icb_rsp_leftover_rdata_nxt = o_icb_rsp_rdata[Y_W-1:0];
  wire [Y_W-1:0] icb_rsp_leftover_rdata_r;
e603_subsys_gnrl_dffl  #(Y_W) icb_rsp_leftover_rdata_dffl (icb_rsp_leftover_ena, icb_rsp_leftover_rdata_nxt, icb_rsp_leftover_rdata_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_err_nxt = o_icb_rsp_err;
  wire icb_rsp_leftover_err_r;
e603_subsys_gnrl_dffl  #(1) icb_rsp_leftover_err_dffl (icb_rsp_leftover_ena, icb_rsp_leftover_err_nxt, icb_rsp_leftover_err_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_excl_ok_nxt = o_icb_rsp_excl_ok;
  wire icb_rsp_leftover_excl_ok_r;
e603_subsys_gnrl_dffl  #(1) icb_rsp_leftover_excl_ok_dffl                   (icb_rsp_leftover_ena, icb_rsp_leftover_excl_ok_nxt, icb_rsp_leftover_excl_ok_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_rsp_leftover_vld = icb_2nd_rsp_valid_r;
  wire i_icb_rsp_valid_cond = (icb_rsp_size_dw ? icb_2nd_rsp_valid_r : 1'b1)
                            ;
  wire o_icb_rsp_ready_byp = (icb_rsp_size_dw & (~icb_2nd_rsp_valid_r))
                             ;
  wire w2n_fifo_o_valid_real = w2n_has_ooo_id_buf ? w2n_fifo_o_match : w2n_fifo_o_valid;
  assign i_icb_rsp_valid =  i_icb_rsp_valid_cond & o_icb_rsp_valid & w2n_fifo_o_valid_real;
  assign i_icb_rsp_rdata = icb_rsp_leftover_vld ? {o_icb_rsp_rdata, icb_rsp_leftover_rdata_r} :
                           icb_rsp_addr_2       ? {o_icb_rsp_rdata, {Y_W{1'b0}}}              :
                                                  {{Y_W{1'b0}}, o_icb_rsp_rdata}
                                                ;
  assign o_icb_rsp_ready = (o_icb_rsp_ready_byp ? 1'b1 : i_icb_rsp_ready) & w2n_fifo_o_valid_real;
  assign i_icb_rsp_err_pre   = icb_rsp_leftover_vld ? (|{icb_rsp_leftover_err_r, o_icb_rsp_err
                                                          }) : 
                                                             (|{
                                                              o_icb_rsp_err
                                                              });
  assign i_icb_rsp_excl_ok_pre = icb_rsp_leftover_vld ? |{icb_rsp_leftover_excl_ok_r, o_icb_rsp_excl_ok} : o_icb_rsp_excl_ok;
  assign i_icb_rsp_usr   = o_icb_rsp_usr;
  generate
    if(SUPPORT_W2N_ID_OOO == 1) begin: rsp_id_ooo_is1
  assign i_icb_rsp_id   = o_icb_rsp_id;
  assign i_icb_rsp_last = icb_rsp_fixed_cvt ? icb_rsp_last : o_icb_rsp_last;
    end
    else begin: rsp_id_ooo_is0
    end
  endgenerate
endmodule
`include "global.v"
module e603_subsys_ficbw2n_gnrl_ooo_id_buf # (
  parameter IDW   = 32,
  parameter DP   = 8,
  parameter DP_PTR_W = 4,
  parameter DW   = 32
) (
  input           i_vld, 
  output          i_rdy, 
  input [IDW-1:0] i_id, 
  input  [DW-1:0] i_dat,
  output          o_vld, 
  output          o_match, 
  input           o_rdy, 
  output [DW-1:0] o_dat,
  input [IDW-1:0] o_id,  
  input           clk,
  input           rst_n
);
genvar i;
integer j;
    wire [DW-1:0] fifo_rf_r [DP-1:0];
    wire [IDW-1:0] fifo_id_r  [DP-1:0];
    wire [DP-1:0]  fifo_vld_set;
    wire [DP-1:0]  fifo_vld_clr;
    wire [DP-1:0]  fifo_vld_ena;
    wire [DP-1:0]  fifo_vld_nxt;
    wire [DP-1:0]  fifo_vld_r;
    wire [DP-1:0]  fifo_dep_set;
    wire [DP-1:0]  fifo_dep_clr;
    wire [DP-1:0]  fifo_dep_ena;
    wire [DP-1:0]  fifo_dep_nxt;
    wire [DP-1:0]  fifo_dep_r;
    wire [DP-1:0]  fifo_last_set;
    wire [DP-1:0]  fifo_last_clr;
    wire [DP-1:0]  fifo_last_ena;
    wire [DP-1:0]  fifo_last_nxt;
    wire [DP-1:0]  fifo_last_r;
    wire [DP_PTR_W-1:0] fifo_dep_entid_r [DP-1:0];
    wire [DP-1:0] fifo_rf_ena;
    wire wen = i_vld & i_rdy;
    wire ren = o_vld & o_rdy;
    wire [DP-1:0] rptr_vec_r;
    wire [DP-1:0] wptr_vec_r;
    wire [DP-1:0] i_id_match_id;
    wire [DP-1:0] i_id_match_id_noclr;
    wire [DP-1:0] i_id_match_id_last;
    reg [DP_PTR_W-1:0] i_id_match_id_entid;
  generate 
    for (i=0; i<DP; i=i+1) begin:gen_wptr_vec
      if(i == 0) begin: i_is_0
          assign wptr_vec_r[i] = (~fifo_vld_r[i]);
      end
      else begin: i_is_not0
          assign wptr_vec_r[i] = (~fifo_vld_r[i]) & (&fifo_vld_r[i-1:0]);
      end
      assign rptr_vec_r[i] = (fifo_vld_r[i] & (o_id == fifo_id_r[i]) & (~fifo_dep_r[i]));
      assign i_id_match_id[i] = (fifo_vld_r[i] & (i_id == fifo_id_r[i]));
      assign i_id_match_id_noclr[i] = i_id_match_id[i] & (~fifo_vld_clr[i]) ;
      assign i_id_match_id_last[i]  = i_id_match_id[i] & fifo_last_r[i] ;
    end
  endgenerate
      assign i_rdy = |(~fifo_vld_r);
  generate 
    for (i=0; i<DP; i=i+1) begin:gen_fifo_rf
      assign fifo_rf_ena[i] = wen & wptr_vec_r[i];
e603_subsys_gnrl_dfflr  #(DW) fifo_rf_dffl (fifo_rf_ena[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(IDW) fifo_id_dffl (fifo_rf_ena[i], i_id , fifo_id_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      assign fifo_vld_set[i] = fifo_rf_ena[i];
      assign fifo_vld_clr[i] = ren & rptr_vec_r[i];
      assign fifo_vld_ena[i] = fifo_vld_set[i] | fifo_vld_clr[i] ;
      assign fifo_vld_nxt[i] = fifo_vld_set[i];
e603_subsys_gnrl_dfflr #(1)  fifo_vld_dfflr (fifo_vld_ena[i], fifo_vld_nxt[i], fifo_vld_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      assign fifo_dep_set[i] = fifo_vld_set[i] & 
                                  (|i_id_match_id_noclr);
// spyglass disable_block ImproperRangeIndex-ML
// SMD: Index fifo_dep_entid_r of width is larger than the width required for the max value of the signal fifo_vld_clr
// SJ:  This is not cared
      assign fifo_dep_clr[i] = fifo_vld_clr[i] | (fifo_dep_r[i] & fifo_vld_clr[fifo_dep_entid_r[i]]);
// spyglass enable_block ImproperRangeIndex-ML
      assign fifo_dep_ena[i] = fifo_dep_set[i] | fifo_dep_clr[i] ;
      assign fifo_dep_nxt[i] = fifo_dep_set[i];
e603_subsys_gnrl_dfflr #(1)  fifo_dep_dffl (fifo_dep_ena[i], fifo_dep_nxt[i], fifo_dep_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      assign fifo_last_set[i] = fifo_vld_set[i]; 
      assign fifo_last_clr[i] = fifo_vld_clr[i] | (fifo_last_r[i] & wen & i_id_match_id[i]);
      assign fifo_last_ena[i] = fifo_last_set[i] | fifo_last_clr[i] ;
      assign fifo_last_nxt[i] = fifo_last_set[i];
e603_subsys_gnrl_dfflr #(1)  fifo_last_dffl (fifo_last_ena[i], fifo_last_nxt[i], fifo_last_r[i], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(DP_PTR_W)              fifo_dep_entid_dffl (fifo_dep_set[i], i_id_match_id_entid, fifo_dep_entid_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
  endgenerate
    always @*
        begin : fifo_dep_entid_nxt_PROC
          i_id_match_id_entid = {DP_PTR_W{1'b0}};
          for(j=0; j<DP; j=j+1) begin
// spyglass disable_block W216
// SMD: Inappropriate range select for int_part_sel variable
// SJ:  Here is not a real issue
            i_id_match_id_entid = i_id_match_id_entid | ({DP_PTR_W{i_id_match_id_last[j]}} & j[DP_PTR_W-1:0]);
// spyglass enable_block W216
          end
        end
    wire [DW-1:0] mux_rdat;
    reg [DW-1:0] mux_rdat_t;
        always @*
        begin : rd_port_PROC
          mux_rdat_t = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_t = mux_rdat_t | ({DW{rptr_vec_r[j]}} & fifo_rf_r[j]);
          end
        end
    assign mux_rdat = mux_rdat_t;
        assign o_dat = mux_rdat;
    assign o_vld = |fifo_vld_r;
    assign o_match = |rptr_vec_r;
endmodule 
module e603_subsys_gnrl_ficb_ww2nn_id # (
    parameter ID_W = 4,
    parameter FIFO_OUTS_CNT_W = 3,
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 0,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 128,
  parameter Y_W = 32
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [ID_W-1:0] i_icb_cmd_id,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W/2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W/16-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [ID_W-1:0]  dw_icb_cmd_id;
  wire [O_AXLEN_W-1:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W/2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
  wire [ID_W-1:0]  dw_icb_rsp_id;
  wire             dw_icb_rsp_last;
  e603_subsys_gnrl_ficb_w2n_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W/2 )
  ) u_ficb_x2x_div2 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id       (i_icb_cmd_id    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id       (i_icb_rsp_id    ),
    .i_icb_rsp_last       (i_icb_rsp_last    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_id       (dw_icb_cmd_id     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .o_icb_rsp_id       (dw_icb_rsp_id     ),
    .o_icb_rsp_last       (dw_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_w2n_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W/2),
    .Y_W(Y_W )
  ) u_ficb_x_div2_to_y (
    .i_icb_cmd_sel       (dw_icb_cmd_sel    ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_id       (dw_icb_cmd_id    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .i_icb_rsp_id       (dw_icb_rsp_id    ),
    .i_icb_rsp_last       (dw_icb_rsp_last    ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id       (o_icb_cmd_id     ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id       (o_icb_rsp_id     ),
    .o_icb_rsp_last       (o_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_www2nnn_id # (
    parameter ID_W = 4,
    parameter FIFO_OUTS_CNT_W = 3,
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 0,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 256,
  parameter Y_W = 32
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [ID_W-1:0] i_icb_cmd_id,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  wire               dw_icb_cmd_sel;
  wire               dw_icb_cmd_valid;
  wire               dw_icb_cmd_ready;
  wire               dw_icb_cmd_read;
  wire [AW-1:0]      dw_icb_cmd_addr;
  wire [X_W/2-1:0]      dw_icb_cmd_wdata;
  wire [(X_W/16-1):0]  dw_icb_cmd_wmask;
  wire               dw_icb_cmd_lock;
  wire               dw_icb_cmd_excl;
  wire [2:0]         dw_icb_cmd_size;
  wire [1:0]         dw_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw_icb_cmd_usr;
  wire [ID_W-1:0]  dw_icb_cmd_id;
  wire [O_AXLEN_W-1:0]         dw_icb_cmd_xlen;
  wire [1:0]         dw_icb_cmd_xburst;
  wire [1:0]         dw_icb_cmd_modes;
  wire               dw_icb_cmd_dmode;
  wire [2:0]         dw_icb_cmd_attri;
  wire               dw_icb_rsp_valid;
  wire               dw_icb_rsp_ready;
  wire               dw_icb_rsp_err;
  wire               dw_icb_rsp_excl_ok;
  wire [X_W/2-1:0]      dw_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw_icb_rsp_usr;
  wire [ID_W-1:0]  dw_icb_rsp_id;
  wire             dw_icb_rsp_last;
 wire                dw2_icb_cmd_sel;
  wire               dw2_icb_cmd_valid;
  wire               dw2_icb_cmd_ready;
  wire               dw2_icb_cmd_read;
  wire [AW-1:0]      dw2_icb_cmd_addr;
  wire [X_W/4-1:0]   dw2_icb_cmd_wdata;
  wire [(X_W/32-1):0]dw2_icb_cmd_wmask;
  wire               dw2_icb_cmd_lock;
  wire               dw2_icb_cmd_excl;
  wire [2:0]         dw2_icb_cmd_size;
  wire [1:0]         dw2_icb_cmd_beat;
  wire [CMD_UW-1:0]  dw2_icb_cmd_usr;
  wire [ID_W-1:0]  dw2_icb_cmd_id;
  wire [O_AXLEN_W-1:0]         dw2_icb_cmd_xlen;
  wire [1:0]         dw2_icb_cmd_xburst;
  wire [1:0]         dw2_icb_cmd_modes;
  wire               dw2_icb_cmd_dmode;
  wire [2:0]         dw2_icb_cmd_attri;
  wire               dw2_icb_rsp_valid;
  wire               dw2_icb_rsp_ready;
  wire               dw2_icb_rsp_err;
  wire               dw2_icb_rsp_excl_ok;
  wire [X_W/4-1:0]   dw2_icb_rsp_rdata;
  wire [RSP_UW-1:0]  dw2_icb_rsp_usr;
  wire [ID_W-1:0]  dw2_icb_rsp_id;
  wire             dw2_icb_rsp_last;
  e603_subsys_gnrl_ficb_w2n_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(X_W/2 )
  ) u_ficb_x2x_div2 (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id       (i_icb_cmd_id    ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id       (i_icb_rsp_id    ),
    .i_icb_rsp_last       (i_icb_rsp_last    ),
    .o_icb_cmd_sel       (dw_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw_icb_cmd_usr     ),
    .o_icb_cmd_id       (dw_icb_cmd_id     ),
    .o_icb_cmd_xlen      (dw_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw_icb_rsp_usr     ),
    .o_icb_rsp_id       (dw_icb_rsp_id     ),
    .o_icb_rsp_last       (dw_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_w2n_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W/2),
    .Y_W(X_W/4)
  ) u_ficb_x_div2_to_x_div4 (
    .i_icb_cmd_sel       (dw_icb_cmd_sel    ),
    .i_icb_cmd_valid     (dw_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw_icb_cmd_usr    ),
    .i_icb_cmd_id       (dw_icb_cmd_id    ),
    .i_icb_cmd_xlen      (dw_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw_icb_rsp_usr    ),
    .i_icb_rsp_id       (dw_icb_rsp_id    ),
    .i_icb_rsp_last       (dw_icb_rsp_last    ),
    .o_icb_cmd_sel       (dw2_icb_cmd_sel     ),
    .o_icb_cmd_valid     (dw2_icb_cmd_valid   ),
    .o_icb_cmd_ready     (dw2_icb_cmd_ready   ),
    .o_icb_cmd_read      (dw2_icb_cmd_read    ),
    .o_icb_cmd_addr      (dw2_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (dw2_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (dw2_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (dw2_icb_cmd_lock    ),
    .o_icb_cmd_excl      (dw2_icb_cmd_excl    ),
    .o_icb_cmd_size      (dw2_icb_cmd_size    ),
    .o_icb_cmd_beat      (dw2_icb_cmd_beat    ),
    .o_icb_cmd_usr       (dw2_icb_cmd_usr     ),
    .o_icb_cmd_id       (dw2_icb_cmd_id     ),
    .o_icb_cmd_xlen      (dw2_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (dw2_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (dw2_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (dw2_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (dw2_icb_cmd_attri   ),
    .o_icb_rsp_valid     (dw2_icb_rsp_valid   ),
    .o_icb_rsp_ready     (dw2_icb_rsp_ready   ),
    .o_icb_rsp_err       (dw2_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (dw2_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (dw2_icb_rsp_usr     ),
    .o_icb_rsp_id       (dw2_icb_rsp_id     ),
    .o_icb_rsp_last       (dw2_icb_rsp_last     ),
    .clk  (clk),
    .rst_n(rst_n)
  );
  e603_subsys_gnrl_ficb_w2n_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W/4),
    .Y_W(Y_W)
  ) u_ficb_x_div4_to_y (
    .i_icb_cmd_sel       (dw2_icb_cmd_sel    ),
    .i_icb_cmd_valid     (dw2_icb_cmd_valid  ),
    .i_icb_cmd_ready     (dw2_icb_cmd_ready  ),
    .i_icb_cmd_read      (dw2_icb_cmd_read   ),
    .i_icb_cmd_addr      (dw2_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (dw2_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (dw2_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (dw2_icb_cmd_lock   ),
    .i_icb_cmd_excl      (dw2_icb_cmd_excl   ),
    .i_icb_cmd_size      (dw2_icb_cmd_size   ),
    .i_icb_cmd_beat      (dw2_icb_cmd_beat   ),
    .i_icb_cmd_usr       (dw2_icb_cmd_usr    ),
    .i_icb_cmd_id        (dw2_icb_cmd_id     ),
    .i_icb_cmd_xlen      (dw2_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (dw2_icb_cmd_xburst ),
    .i_icb_cmd_modes     (dw2_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (dw2_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (dw2_icb_cmd_attri  ),
    .i_icb_rsp_valid     (dw2_icb_rsp_valid  ),
    .i_icb_rsp_ready     (dw2_icb_rsp_ready  ),
    .i_icb_rsp_err       (dw2_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (dw2_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (dw2_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (dw2_icb_rsp_usr    ),
    .i_icb_rsp_id        (dw2_icb_rsp_id     ),
    .i_icb_rsp_last        (dw2_icb_rsp_last     ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id        (o_icb_cmd_id      ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id        (o_icb_rsp_id      ),
    .o_icb_rsp_last        (o_icb_rsp_last      ),
    .clk  (clk),
    .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb_wconv_id # (
    parameter ID_W = 4,
    parameter FIFO_OUTS_CNT_W = 3,
    parameter SUPPORT_W2N_ID_OOO = 0,
  parameter O_AXLEN_EXTEND = 0, 
  parameter O_AXLEN_W = 8, 
  parameter PAYLOAD_NORST = 0,
  parameter ZEROCYC_RSP = 0,
  parameter AW = 64,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1,
  parameter RSP_CHECK_CMD_OUTS = 0,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 64
) (
  input              i_icb_cmd_sel,
  input              i_icb_cmd_valid,
  output             i_icb_cmd_ready,
  input              i_icb_cmd_read,
  input  [AW-1:0]    i_icb_cmd_addr,
  input  [X_W-1:0]   i_icb_cmd_wdata,
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [O_AXLEN_W-1:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  input  [ID_W-1:0] i_icb_cmd_id,
  output             i_icb_rsp_valid,
  input              i_icb_rsp_ready,
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel,
  output             o_icb_cmd_valid,
  input              o_icb_cmd_ready,
  output             o_icb_cmd_read,
  output [AW-1:0]    o_icb_cmd_addr,
  output [Y_W-1:0]   o_icb_cmd_wdata,
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [O_AXLEN_W-1:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid,
  output             o_icb_rsp_ready,
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata,
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  generate
    if(X_W == Y_W) begin: x_is_y_gen
    wire rspid_fifo_i_ready;
    wire rspid_fifo_o_valid;
        if(RSP_CHECK_CMD_OUTS == 1) begin: rsp_fifo_gen
    wire rspid_fifo_i_push = o_icb_cmd_valid & o_icb_cmd_ready
                           ;
    wire rspid_fifo_o_pop  = o_icb_rsp_valid & o_icb_rsp_ready
                           ;
    e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT(1'b1),
        .CUT_READY (FIFO_CUT_READY),
        .DP  (FIFO_OUTS_NUM+1),
        .DW  (1)
      ) u_e603_subsys_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_push ),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(1'b0 ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_pop),
        .o_dat(),
        .clk  (clk),
        .rst_n(rst_n)
      );
        end
        else begin : no_rsp_fifo_gen
    assign rspid_fifo_i_ready = 1'b1;
    assign rspid_fifo_o_valid = 1'b1;
        end
        assign o_icb_cmd_sel   = i_icb_cmd_sel;
        assign i_icb_cmd_ready = rspid_fifo_i_ready & o_icb_cmd_ready;
        assign o_icb_cmd_valid = rspid_fifo_i_ready & i_icb_cmd_valid;
        assign o_icb_cmd_read  = i_icb_cmd_read ;
        assign o_icb_cmd_addr  = i_icb_cmd_addr ;
        assign o_icb_cmd_wdata = i_icb_cmd_wdata;
        assign o_icb_cmd_wmask = i_icb_cmd_wmask;
        assign o_icb_cmd_beat  = i_icb_cmd_beat ;
        assign o_icb_cmd_lock  = i_icb_cmd_lock ;
        assign o_icb_cmd_excl  = i_icb_cmd_excl ;
        assign o_icb_cmd_size  = i_icb_cmd_size ;
        assign o_icb_cmd_usr   = i_icb_cmd_usr  ;
        assign o_icb_cmd_id    = i_icb_cmd_id   ;
        assign o_icb_cmd_xlen  = i_icb_cmd_xlen  ;
        assign o_icb_cmd_xburst= i_icb_cmd_xburst;
        assign o_icb_cmd_modes = i_icb_cmd_modes ;
        assign o_icb_cmd_dmode = i_icb_cmd_dmode ;
        assign o_icb_cmd_attri = i_icb_cmd_attri ;
        assign o_icb_rsp_ready     = rspid_fifo_o_valid & i_icb_rsp_ready;
        assign i_icb_rsp_valid     = rspid_fifo_o_valid & o_icb_rsp_valid;
        assign i_icb_rsp_err       = o_icb_rsp_err  ;
        assign i_icb_rsp_excl_ok   = o_icb_rsp_excl_ok  ;
        assign i_icb_rsp_rdata     = o_icb_rsp_rdata;
        assign i_icb_rsp_usr       = o_icb_rsp_usr;
        assign i_icb_rsp_id        = o_icb_rsp_id ;
        assign i_icb_rsp_last        = o_icb_rsp_last ;
    end
    if(    ((Y_W ==  64) && (X_W ==  32)) 
        || ((Y_W == 128) && (X_W ==  64))
        || ((Y_W == 256) && (X_W == 128))
        || ((Y_W == 512) && (X_W == 256))
        || ((Y_W == 1024) && (X_W == 512))
        || ((Y_W == 2048) && (X_W == 1024))
        ) begin:n2w_gen
  e603_subsys_gnrl_ficb_n2w_id # (
    .ID_W(ID_W),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_n2w (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id        (i_icb_cmd_id     ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id        (i_icb_rsp_id     ),
    .i_icb_rsp_last        (i_icb_rsp_last     ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id        (o_icb_cmd_id      ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id        (o_icb_rsp_id      ),
    .o_icb_rsp_last        (o_icb_rsp_last      ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((Y_W == 128) && (X_W == 32))
      || ((Y_W == 256) && (X_W == 64))
      || ((Y_W == 512) && (X_W == 128))
      || ((Y_W == 1024) && (X_W == 256))
      || ((Y_W == 2048) && (X_W == 512))
        ) begin:nn2ww_gen
  e603_subsys_gnrl_ficb_nn2ww_id # (
    .ID_W(ID_W),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_nn2ww (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id        (i_icb_cmd_id     ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id        (i_icb_rsp_id     ),
    .i_icb_rsp_last        (i_icb_rsp_last     ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id        (o_icb_cmd_id      ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id        (o_icb_rsp_id      ),
    .o_icb_rsp_last        (o_icb_rsp_last      ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((Y_W == 256) && (X_W == 32))
      || ((Y_W == 512) && (X_W == 64))
      || ((Y_W == 1024) && (X_W == 128))
      || ((Y_W == 2048) && (X_W == 256))
        ) begin:nnn2www_gen
  e603_subsys_gnrl_ficb_nnn2www_id # (
    .ID_W(ID_W),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_nnn2www (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id        (i_icb_cmd_id     ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id        (i_icb_rsp_id     ),
    .i_icb_rsp_last        (i_icb_rsp_last     ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id        (o_icb_cmd_id      ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id        (o_icb_rsp_id      ),
    .o_icb_rsp_last        (o_icb_rsp_last      ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(    ((X_W ==  64) && (Y_W ==  32)) 
        || ((X_W == 128) && (Y_W ==  64))
        || ((X_W == 256) && (Y_W == 128))
        || ((X_W == 512) && (Y_W == 256))
        || ((X_W == 1024) && (Y_W == 512))
        ) begin:w2n_gen
  e603_subsys_gnrl_ficb_w2n_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_w2n (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id        (i_icb_cmd_id     ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id        (i_icb_rsp_id     ),
    .i_icb_rsp_last        (i_icb_rsp_last     ),
    .o_icb_cmd_sel       (o_icb_cmd_sel     ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id        (o_icb_cmd_id      ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id        (o_icb_rsp_id      ),
    .o_icb_rsp_last        (o_icb_rsp_last      ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((X_W == 128) && (Y_W == 32))
      || ((X_W == 256) && (Y_W == 64))
      || ((X_W == 512) && (Y_W == 128))
      || ((X_W == 1024) && (Y_W == 256))
        ) begin:ww2nn
  e603_subsys_gnrl_ficb_ww2nn_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_ww2nn (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id        (i_icb_cmd_id     ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id        (i_icb_rsp_id     ),
    .i_icb_rsp_last        (i_icb_rsp_last     ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id        (o_icb_cmd_id      ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id        (o_icb_rsp_id      ),
    .o_icb_rsp_last        (o_icb_rsp_last      ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
    if(
         ((X_W == 256) && (Y_W == 32))
      || ((X_W == 512) && (Y_W == 64))
      || ((X_W == 1024) && (Y_W == 128))
        ) begin:www2nnn
  e603_subsys_gnrl_ficb_www2nnn_id # (
    .ID_W(ID_W),
    .FIFO_OUTS_CNT_W(FIFO_OUTS_CNT_W),
    .SUPPORT_W2N_ID_OOO(SUPPORT_W2N_ID_OOO),
    .ZEROCYC_RSP   (ZEROCYC_RSP   ),
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .AW            (AW            ),
    .CMD_UW        (CMD_UW        ),
    .RSP_UW        (RSP_UW        ),
    .FIFO_OUTS_NUM (FIFO_OUTS_NUM ),
    .FIFO_CUT_READY(FIFO_CUT_READY),
    .X_W(X_W),
    .Y_W(Y_W )
  ) u_ficb_www2nnn (
    .i_icb_cmd_sel       (i_icb_cmd_sel    ),
    .i_icb_cmd_valid     (i_icb_cmd_valid  ),
    .i_icb_cmd_ready     (i_icb_cmd_ready  ),
    .i_icb_cmd_read      (i_icb_cmd_read   ),
    .i_icb_cmd_addr      (i_icb_cmd_addr   ),
    .i_icb_cmd_wdata     (i_icb_cmd_wdata  ),
    .i_icb_cmd_wmask     (i_icb_cmd_wmask  ),
    .i_icb_cmd_lock      (i_icb_cmd_lock   ),
    .i_icb_cmd_excl      (i_icb_cmd_excl   ),
    .i_icb_cmd_size      (i_icb_cmd_size   ),
    .i_icb_cmd_beat      (i_icb_cmd_beat   ),
    .i_icb_cmd_usr       (i_icb_cmd_usr    ),
    .i_icb_cmd_id        (i_icb_cmd_id     ),
    .i_icb_cmd_xlen      (i_icb_cmd_xlen   ),
    .i_icb_cmd_xburst    (i_icb_cmd_xburst ),
    .i_icb_cmd_modes     (i_icb_cmd_modes  ),
    .i_icb_cmd_dmode     (i_icb_cmd_dmode  ),
    .i_icb_cmd_attri     (i_icb_cmd_attri  ),
    .i_icb_rsp_valid     (i_icb_rsp_valid  ),
    .i_icb_rsp_ready     (i_icb_rsp_ready  ),
    .i_icb_rsp_err       (i_icb_rsp_err    ),
    .i_icb_rsp_excl_ok   (i_icb_rsp_excl_ok),
    .i_icb_rsp_rdata     (i_icb_rsp_rdata  ),
    .i_icb_rsp_usr       (i_icb_rsp_usr    ),
    .i_icb_rsp_id        (i_icb_rsp_id     ),
    .i_icb_rsp_last        (i_icb_rsp_last     ),
    .o_icb_cmd_sel       (o_icb_cmd_sel   ),
    .o_icb_cmd_valid     (o_icb_cmd_valid   ),
    .o_icb_cmd_ready     (o_icb_cmd_ready   ),
    .o_icb_cmd_read      (o_icb_cmd_read    ),
    .o_icb_cmd_addr      (o_icb_cmd_addr    ),
    .o_icb_cmd_wdata     (o_icb_cmd_wdata   ),
    .o_icb_cmd_wmask     (o_icb_cmd_wmask   ),
    .o_icb_cmd_lock      (o_icb_cmd_lock    ),
    .o_icb_cmd_excl      (o_icb_cmd_excl    ),
    .o_icb_cmd_size      (o_icb_cmd_size    ),
    .o_icb_cmd_beat      (o_icb_cmd_beat    ),
    .o_icb_cmd_usr       (o_icb_cmd_usr     ),
    .o_icb_cmd_id        (o_icb_cmd_id      ),
    .o_icb_cmd_xlen      (o_icb_cmd_xlen    ),
    .o_icb_cmd_xburst    (o_icb_cmd_xburst  ),
    .o_icb_cmd_modes     (o_icb_cmd_modes   ),
    .o_icb_cmd_dmode     (o_icb_cmd_dmode   ),
    .o_icb_cmd_attri     (o_icb_cmd_attri   ),
    .o_icb_rsp_valid     (o_icb_rsp_valid   ),
    .o_icb_rsp_ready     (o_icb_rsp_ready   ),
    .o_icb_rsp_err       (o_icb_rsp_err     ),
    .o_icb_rsp_excl_ok   (o_icb_rsp_excl_ok ),
    .o_icb_rsp_rdata     (o_icb_rsp_rdata   ),
    .o_icb_rsp_usr       (o_icb_rsp_usr     ),
    .o_icb_rsp_id        (o_icb_rsp_id      ),
    .o_icb_rsp_last        (o_icb_rsp_last      ),
    .clk  (clk),
    .rst_n(rst_n)
  );
    end
  endgenerate
endmodule
module e603_subsys_gnrl_ficb_splt_id
 # (
    parameter ID_W = 4,
  parameter AW = 32,
  parameter DW = 64,
  parameter USE_ALL_READY = 0,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter SPLT_NUM = 4,
  parameter SPLT_PTR_1HOT = 1,
  parameter PAYLOAD_NORST = 0,
  parameter SPLT_PTR_W = 4,
  parameter FIFO_REG_OUT = 0,
  parameter ALLOW_DIFF = 1,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  input  [SPLT_NUM-1:0] i_icb_splt_indic,
  input  [SPLT_NUM-1:0] o_icb_support_oid,
  output splt_active,
  input  clk_en,
  input  i_icb_cmd_sel,
  input  i_icb_cmd_valid,
  output i_icb_cmd_ready,
  input             i_icb_cmd_read,
  input  [AW-1:0]   i_icb_cmd_addr,
  input  [DW-1:0]   i_icb_cmd_wdata,
  input  [DW/8-1:0]   i_icb_cmd_wmask,
  input  [1:0]      i_icb_cmd_beat,
  input             i_icb_cmd_lock,
  input             i_icb_cmd_excl,
  input  [2:0]      i_icb_cmd_size,
  input  [CMD_UW-1:0]i_icb_cmd_usr,
  input [7:0]       i_icb_cmd_xlen,
  input [1:0]       i_icb_cmd_xburst,
  input [1:0]       i_icb_cmd_modes,
  input             i_icb_cmd_dmode,
  input [2:0]       i_icb_cmd_attri,
  input  [ID_W-1:0] i_icb_cmd_id,
  output i_icb_rsp_valid,
  input  i_icb_rsp_ready,
  output i_icb_rsp_err,
  output i_icb_rsp_excl_ok,
  output [DW-1:0] i_icb_rsp_rdata,
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  input  [SPLT_NUM*1-1:0]    o_bus_icb_cmd_ready,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_valid,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_sel,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_read,
  output [SPLT_NUM*AW-1:0]   o_bus_icb_cmd_addr,
  output [SPLT_NUM*DW-1:0]   o_bus_icb_cmd_wdata,
  output [SPLT_NUM*DW/8-1:0]   o_bus_icb_cmd_wmask,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_beat,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_lock,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_excl,
  output [SPLT_NUM*3-1:0]    o_bus_icb_cmd_size,
  output [SPLT_NUM*CMD_UW-1:0]o_bus_icb_cmd_usr,
  output [SPLT_NUM*ID_W-1:0]  o_bus_icb_cmd_id,
  output [SPLT_NUM*8-1:0]    o_bus_icb_cmd_xlen,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_xburst,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_modes,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_dmode,
  output [SPLT_NUM*3-1:0]    o_bus_icb_cmd_attri,
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_valid,
  output [SPLT_NUM*1-1:0]  o_bus_icb_rsp_ready,
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_err,
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_excl_ok,
  input  [SPLT_NUM*DW-1:0] o_bus_icb_rsp_rdata,
  input  [SPLT_NUM*RSP_UW-1:0] o_bus_icb_rsp_usr,
  input  [SPLT_NUM*ID_W-1:0] o_bus_icb_rsp_id,
  input  [SPLT_NUM     -1:0] o_bus_icb_rsp_last,
  input  clk,
  input  rst_n
  );
  wire [SPLT_NUM-1:0] i_icb_splt_indic_real;
    wire i_icb_cmd_hsked = i_icb_cmd_valid & i_icb_cmd_ready;
    assign i_icb_splt_indic_real = i_icb_splt_indic;
  localparam SPLT_FIFO_DW = (SPLT_PTR_W + ID_W + 1) 
                       ;
  wire rspid_fifo_empty;
generate 
  if(SPLT_NUM == 1) begin:gen_splt_num_eq_1
    assign i_icb_cmd_ready     = o_bus_icb_cmd_ready;
    assign o_bus_icb_cmd_sel   = i_icb_cmd_sel;
    assign o_bus_icb_cmd_valid = i_icb_cmd_valid;
    assign o_bus_icb_cmd_read  = i_icb_cmd_read ;
    assign o_bus_icb_cmd_addr  = i_icb_cmd_addr ;
    assign o_bus_icb_cmd_wdata = i_icb_cmd_wdata;
    assign o_bus_icb_cmd_wmask = i_icb_cmd_wmask;
    assign o_bus_icb_cmd_beat  = i_icb_cmd_beat ;
    assign o_bus_icb_cmd_lock  = i_icb_cmd_lock ;
    assign o_bus_icb_cmd_excl  = i_icb_cmd_excl ;
    assign o_bus_icb_cmd_size  = i_icb_cmd_size ;
    assign o_bus_icb_cmd_usr   = i_icb_cmd_usr  ;
    assign o_bus_icb_cmd_id    = i_icb_cmd_id  ;
    assign o_bus_icb_cmd_xlen  = i_icb_cmd_xlen  ;
    assign o_bus_icb_cmd_xburst= i_icb_cmd_xburst;
    assign o_bus_icb_cmd_modes = i_icb_cmd_modes ;
    assign o_bus_icb_cmd_dmode = i_icb_cmd_dmode ;
    assign o_bus_icb_cmd_attri = i_icb_cmd_attri ;
    assign rspid_fifo_empty    = 1'b1;
    assign o_bus_icb_rsp_ready = i_icb_rsp_ready;
    assign i_icb_rsp_valid     = o_bus_icb_rsp_valid;
    assign i_icb_rsp_err       = o_bus_icb_rsp_err  ;
    assign i_icb_rsp_excl_ok   = o_bus_icb_rsp_excl_ok  ;
    assign i_icb_rsp_rdata     = o_bus_icb_rsp_rdata;
    assign i_icb_rsp_usr       = o_bus_icb_rsp_usr;
    assign i_icb_rsp_id        = o_bus_icb_rsp_id ;
    assign i_icb_rsp_last        = o_bus_icb_rsp_last ;
  end
  else begin:gen_splt_num_gt_1
    genvar i;
    genvar ii;
    integer j;
    wire [SPLT_NUM-1:0] o_icb_cmd_sel;
    wire [SPLT_NUM-1:0] o_icb_cmd_valid;
    wire [SPLT_NUM-1:0] o_icb_cmd_ready;
    wire            o_icb_cmd_read [SPLT_NUM-1:0];
    wire [AW-1:0]   o_icb_cmd_addr [SPLT_NUM-1:0];
    wire [DW-1:0]   o_icb_cmd_wdata[SPLT_NUM-1:0];
    wire [DW/8-1:0]   o_icb_cmd_wmask[SPLT_NUM-1:0];
    wire [1:0]      o_icb_cmd_beat [SPLT_NUM-1:0];
    wire            o_icb_cmd_lock [SPLT_NUM-1:0];
    wire            o_icb_cmd_excl [SPLT_NUM-1:0];
    wire [2:0]      o_icb_cmd_size [SPLT_NUM-1:0];
    wire [CMD_UW-1:0]o_icb_cmd_usr  [SPLT_NUM-1:0];
    wire [7:0]      o_icb_cmd_xlen  [SPLT_NUM-1:0];
    wire [1:0]      o_icb_cmd_xburst[SPLT_NUM-1:0];
    wire [1:0]      o_icb_cmd_modes [SPLT_NUM-1:0];
    wire            o_icb_cmd_dmode [SPLT_NUM-1:0];
    wire [2:0]      o_icb_cmd_attri [SPLT_NUM-1:0];
    wire [ID_W-1:0] o_icb_cmd_id [SPLT_NUM-1:0];
    wire [SPLT_NUM-1:0] o_icb_rsp_valid;
    wire [SPLT_NUM-1:0] o_icb_rsp_ready;
    wire [SPLT_NUM-1:0] o_icb_rsp_err  ;
    wire [SPLT_NUM-1:0] o_icb_rsp_excl_ok  ;
    wire [DW-1:0] o_icb_rsp_rdata  [SPLT_NUM-1:0];
    wire [RSP_UW-1:0] o_icb_rsp_usr [SPLT_NUM-1:0];
    wire [ID_W-1:0] o_icb_rsp_id [SPLT_NUM-1:0];
    wire [SPLT_NUM-1:0] o_icb_rsp_last;
    wire [SPLT_NUM-1:0] o_icb_cmd_ready_excpt_this [SPLT_NUM-1:0];
    wire sel_o_icb_cmd_ready;
    wire rspid_fifo_bypass;
    wire rspid_fifo_wen;
    wire rspid_fifo_ren;
    wire [SPLT_PTR_W-1:0] o_icb_rsp_port_id;
    wire rspid_fifo_i_valid;
    wire rspid_fifo_o_valid;
    wire rspid_fifo_o_valid_real;
    wire rspid_fifo_i_ready;
    wire rspid_fifo_i_ready_real;
    wire rspid_fifo_o_ready;
    wire [SPLT_FIFO_DW-1:0] rspid_fifo_rdat;
    wire [SPLT_FIFO_DW-1:0] rspid_fifo_rdat_real;
    wire [SPLT_FIFO_DW-1:0] rspid_fifo_wdat;
    wire rspid_fifo_full;
    reg [SPLT_PTR_W-1:0] i_splt_indic_id;
    wire i_icb_cmd_ready_pre;
    wire i_icb_cmd_valid_pre;
    wire i_icb_cmd_sel_pre;
    wire cmd_diff_branch_t[SPLT_NUM-1:0];
    wire i_icb_cmd_valid_pre2[SPLT_NUM-1:0];
    wire i_icb_cmd_sel_pre2[SPLT_NUM-1:0];
    wire i_icb_rsp_ready_pre;
    wire i_icb_rsp_valid_pre;
    for(i = 0; i < SPLT_NUM; i = i+1)
    begin:gen_icb_distract
      assign o_icb_cmd_ready[i]                             = o_bus_icb_cmd_ready[(i+1)*1     -1 : (i)*1     ];
      assign o_bus_icb_cmd_sel  [(i+1)*1     -1 : i*1     ] = o_icb_cmd_sel[i];
      assign o_bus_icb_cmd_valid[(i+1)*1     -1 : i*1     ] = o_icb_cmd_valid[i];
      assign o_bus_icb_cmd_read [(i+1)*1     -1 : i*1     ] = o_icb_cmd_read [i];
      assign o_bus_icb_cmd_addr [(i+1)*AW    -1 : i*AW    ] = o_icb_cmd_addr [i];
      assign o_bus_icb_cmd_wdata[(i+1)*DW    -1 : i*DW    ] = o_icb_cmd_wdata[i];
      assign o_bus_icb_cmd_wmask[(i+1)*DW/8    -1 : i*DW/8    ] = o_icb_cmd_wmask[i];
      assign o_bus_icb_cmd_beat [(i+1)*2     -1 : i*2     ] = o_icb_cmd_beat [i];
      assign o_bus_icb_cmd_lock [(i+1)*1     -1 : i*1     ] = o_icb_cmd_lock [i];
      assign o_bus_icb_cmd_excl [(i+1)*1     -1 : i*1     ] = o_icb_cmd_excl [i];
      assign o_bus_icb_cmd_size [(i+1)*3     -1 : i*3     ] = o_icb_cmd_size [i];
      assign o_bus_icb_cmd_usr  [(i+1)*CMD_UW -1 : i*CMD_UW ] = o_icb_cmd_usr  [i];
      assign o_bus_icb_cmd_xlen  [(i+1)*8 -1 : i*8 ] = o_icb_cmd_xlen  [i];
      assign o_bus_icb_cmd_xburst[(i+1)*2 -1 : i*2 ] = o_icb_cmd_xburst[i];
      assign o_bus_icb_cmd_modes [(i+1)*2 -1 : i*2 ] = o_icb_cmd_modes [i];
      assign o_bus_icb_cmd_dmode [(i+1)*1 -1 : i*1 ] = o_icb_cmd_dmode [i];
      assign o_bus_icb_cmd_attri [(i+1)*3 -1 : i*3 ] = o_icb_cmd_attri [i];
      assign o_bus_icb_cmd_id    [(i+1)*ID_W -1 : i*ID_W ] = o_icb_cmd_id    [i];
      assign o_bus_icb_rsp_ready[(i+1)*1-1 :i*1 ] = o_icb_rsp_ready[i];
      assign o_icb_rsp_valid[i]                   = o_bus_icb_rsp_valid[(i+1)*1-1 :i*1 ];
      assign o_icb_rsp_err  [i]                   = o_bus_icb_rsp_err  [(i+1)*1-1 :i*1 ];
      assign o_icb_rsp_excl_ok  [i]               = o_bus_icb_rsp_excl_ok  [(i+1)*1-1 :i*1 ];
      assign o_icb_rsp_rdata[i]                   = o_bus_icb_rsp_rdata[(i+1)*DW-1:i*DW];
      assign o_icb_rsp_usr       [i]              = o_bus_icb_rsp_usr  [(i+1)*RSP_UW-1:i*RSP_UW];
      assign { o_icb_rsp_last[i], 
                 o_icb_rsp_id[i]
                 }              = 
                                o_icb_support_oid[i] ?   
                               {
                                                     o_bus_icb_rsp_last[(i+1)*1-1 :i*1 ],
                                                     o_bus_icb_rsp_id  [(i+1)*ID_W-1:i*ID_W]
                                }
                                                     : {
                                                         rspid_fifo_rdat_real[SPLT_PTR_W+ID_W],
                                                         rspid_fifo_rdat_real[SPLT_PTR_W+ID_W-1:SPLT_PTR_W] 
                                                         } 
                                                         ;
    end
    if(USE_ALL_READY == 1) begin:gen_all_ready
      assign sel_o_icb_cmd_ready = (&o_icb_cmd_ready);
    end
    else begin:gen_non_all_ready
      reg  sel_o_icb_cmd_ready_reg;
      always @ (*) begin : sel_o_icb_cmd_ready_PROC
        sel_o_icb_cmd_ready_reg = 1'b0;
          for(j = 0; j < SPLT_NUM; j = j+1) begin
            sel_o_icb_cmd_ready_reg = sel_o_icb_cmd_ready_reg | (i_icb_splt_indic_real[j] & o_icb_cmd_ready[j]);
          end
      end
      assign sel_o_icb_cmd_ready = sel_o_icb_cmd_ready_reg;
    end
    assign i_icb_cmd_ready_pre = sel_o_icb_cmd_ready;
    if(ALLOW_DIFF == 1) begin:gen_allow_diff
       assign i_icb_cmd_sel_pre       = i_icb_cmd_sel       & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre     = i_icb_cmd_valid     & (~rspid_fifo_full);
          for(i = 0; i < SPLT_NUM; i = i+1) begin:gen_allow_diff_splt_cmd
       assign cmd_diff_branch_t[i] = 1'b0;
       assign i_icb_cmd_sel_pre2  [i] = i_icb_cmd_sel       & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre2[i] = i_icb_cmd_valid     & (~rspid_fifo_full);
          end
       assign i_icb_cmd_ready     = i_icb_cmd_ready_pre & (~rspid_fifo_full);
    end
    else begin:gen_not_allow_diff
       wire cmd_diff_branch = (~rspid_fifo_empty) & (~(rspid_fifo_wdat[SPLT_PTR_W-1:0] == rspid_fifo_rdat_real[SPLT_PTR_W-1:0]));
       assign i_icb_cmd_sel_pre       = i_icb_cmd_sel       & (~cmd_diff_branch) & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre     = i_icb_cmd_valid     & (~cmd_diff_branch) & (~rspid_fifo_full);
        if(SPLT_PTR_1HOT == 1) begin:gen_pre2_ptr_1hot
          for(i = 0; i < SPLT_NUM; i = i+1) begin:gen_not_allow_diff_splt_cmd
       assign cmd_diff_branch_t[i] = (~rspid_fifo_empty) & (~(rspid_fifo_wdat[i] == rspid_fifo_rdat_real[i]));
       assign i_icb_cmd_sel_pre2   [i] = i_icb_cmd_sel       & (~cmd_diff_branch_t[i]) & (~rspid_fifo_full);
       assign i_icb_cmd_valid_pre2 [i] = i_icb_cmd_valid     & (~cmd_diff_branch_t[i]) & (~rspid_fifo_full);
          end
        end
        else begin: gen_pre2_ptr_not_1hot
          for(i = 0; i < SPLT_NUM; i = i+1) begin:gen_not_allow_diff_splt_cmd
       assign cmd_diff_branch_t[i] = 1'b0;
       assign i_icb_cmd_sel_pre2   [i] = i_icb_cmd_sel_pre;
       assign i_icb_cmd_valid_pre2 [i] = i_icb_cmd_valid_pre;
          end
        end
       assign i_icb_cmd_ready     = i_icb_cmd_ready_pre & (~cmd_diff_branch) & (~rspid_fifo_full);
    end
    if(SPLT_PTR_1HOT == 1) begin:gen_ptr_1hot
       always @ (*) begin : i_splt_indic_id_PROC
         i_splt_indic_id = i_icb_splt_indic_real;
       end
    end
    else begin:gen_ptr_not_1hot
       always @ (*) begin : i_splt_indic_id_PROC
         i_splt_indic_id = {SPLT_PTR_W{1'b0}};
         for(j = 0; j < SPLT_NUM; j = j+1) begin
// spyglass disable_block W216
// SMD: Inappropriate range select for int_part_sel variable
// SJ:  Here is not a real issue
           i_splt_indic_id = i_splt_indic_id | ({SPLT_PTR_W{i_icb_splt_indic_real[j]}} & (j[SPLT_PTR_W-1:0]));
// spyglass enable_block W216
         end
       end
    end
 if(ALLOW_DIFF == 1) begin:rspfifo_gen_allow_diff1
    assign rspid_fifo_wen = i_icb_cmd_valid & i_icb_cmd_ready;
    assign rspid_fifo_ren = i_icb_rsp_valid & i_icb_rsp_ready;
 end
 else begin: rspfifo_gen_allow_diff0
    assign rspid_fifo_wen = i_icb_cmd_valid & i_icb_cmd_ready 
                          ;
    assign rspid_fifo_ren = i_icb_rsp_valid & i_icb_rsp_ready 
                          ;
 end
    if(ALLOW_0CYCL_RSP == 1) begin: gen_allow_0rsp
        assign rspid_fifo_bypass = rspid_fifo_empty & rspid_fifo_wen & rspid_fifo_ren;
        assign o_icb_rsp_port_id = rspid_fifo_empty ? rspid_fifo_wdat[SPLT_PTR_W-1:0] : rspid_fifo_rdat_real[SPLT_PTR_W-1:0];
        assign i_icb_rsp_valid     = i_icb_rsp_valid_pre;
        assign i_icb_rsp_ready_pre = i_icb_rsp_ready;
    end
    else begin: gen_no_allow_0rsp
        assign rspid_fifo_bypass = 1'b0;
        assign o_icb_rsp_port_id = rspid_fifo_rdat_real[SPLT_PTR_W-1:0];
        assign i_icb_rsp_valid     = (~rspid_fifo_empty) & i_icb_rsp_valid_pre;
        assign i_icb_rsp_ready_pre = (~rspid_fifo_empty) & i_icb_rsp_ready;
    end
    assign rspid_fifo_i_valid = clk_en & rspid_fifo_wen & (~rspid_fifo_bypass);
    assign rspid_fifo_full    = (~rspid_fifo_i_ready_real);
    assign rspid_fifo_o_ready = clk_en & rspid_fifo_ren & (~rspid_fifo_bypass);
    assign rspid_fifo_empty   = (~rspid_fifo_o_valid_real);
      wire i_icb_cmd_last = i_icb_cmd_beat[1] | (i_icb_cmd_xlen == 8'd0);
      wire i_icb_cmd_fixed = (i_icb_cmd_xburst == 2'b00);
      assign rspid_fifo_wdat   = {
                               i_icb_cmd_last, i_icb_cmd_id,i_splt_indic_id};
    assign rspid_fifo_o_valid_real = rspid_fifo_o_valid;
    assign rspid_fifo_i_ready_real = rspid_fifo_i_ready;
    assign rspid_fifo_rdat_real = rspid_fifo_rdat;
    if(FIFO_OUTS_NUM == 1) begin:gen_fifo_dp_1
      e603_subsys_gnrl_pipe_stage # (
        .CUT_READY (FIFO_CUT_READY),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (1),
        .DW  (SPLT_FIFO_DW)
      ) u_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    else begin: gen_fifo_dp_gt_1
      e603_subsys_gnrl_fifo # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
        .REG_OUT(FIFO_REG_OUT),
        .CUT_READY (FIFO_CUT_READY),
        .DP  (FIFO_OUTS_NUM),
        .DW  (SPLT_FIFO_DW)
      ) u_gnrl_rspid_fifo (
        .i_vld(rspid_fifo_i_valid),
        .i_rdy(rspid_fifo_i_ready),
        .i_dat(rspid_fifo_wdat ),
        .o_vld(rspid_fifo_o_valid),
        .o_rdy(rspid_fifo_o_ready),
        .o_dat(rspid_fifo_rdat ),
        .clk  (clk),
        .rst_n(rst_n)
      );
    end
    for(i = 0; i < SPLT_NUM; i = i+1)
    begin:gen_o_icb_cmd_valid
      for(ii = 0; ii < SPLT_NUM; ii = ii+1)
      begin:gen_o_cmd_ready_excpt_this
         if(i == ii) begin: gen_same_i
           assign o_icb_cmd_ready_excpt_this[i][ii] = 1'b1;
         end
         else begin: gen_no_same_i
           assign o_icb_cmd_ready_excpt_this[i][ii] = o_icb_cmd_ready[ii];
         end
      end
      if(USE_ALL_READY == 1) begin:gen_all_ready
         assign o_icb_cmd_valid[i] = i_icb_splt_indic_real[i] & i_icb_cmd_valid_pre2[i] & (&o_icb_cmd_ready_excpt_this[i]);
         assign o_icb_cmd_sel  [i] = i_icb_splt_indic_real[i] & i_icb_cmd_sel_pre2[i]   & (&o_icb_cmd_ready_excpt_this[i]);
      end
      else begin:gen_non_all_ready
         assign o_icb_cmd_valid[i] = i_icb_splt_indic_real[i] & i_icb_cmd_valid_pre2[i];
         assign o_icb_cmd_sel  [i] = i_icb_splt_indic_real[i] & i_icb_cmd_sel_pre2[i];
      end
      assign o_icb_cmd_lock[i] = i_icb_cmd_lock;
          assign o_icb_cmd_read [i] = i_icb_cmd_read ;
          assign o_icb_cmd_addr [i] = i_icb_cmd_addr ;
          assign o_icb_cmd_wdata[i] = i_icb_cmd_wdata;
          assign o_icb_cmd_wmask[i] = i_icb_cmd_wmask;
          assign o_icb_cmd_excl [i] = i_icb_cmd_excl ;
          assign o_icb_cmd_size [i] = i_icb_cmd_size ;
          assign o_icb_cmd_usr  [i] = i_icb_cmd_usr  ;
          assign o_icb_cmd_xburst[i] = i_icb_cmd_xburst;
          assign o_icb_cmd_modes [i] = i_icb_cmd_modes ;
          assign o_icb_cmd_dmode [i] = i_icb_cmd_dmode ;
          assign o_icb_cmd_attri [i] = i_icb_cmd_attri ;
          assign o_icb_cmd_xlen  [i] = i_icb_cmd_fixed ? (o_icb_support_oid[i] ? i_icb_cmd_xlen : 8'b0) : i_icb_cmd_xlen;
          assign o_icb_cmd_beat  [i] = i_icb_cmd_fixed ? (o_icb_support_oid[i] ? i_icb_cmd_beat : 2'b0) : i_icb_cmd_beat;
          assign o_icb_cmd_id [i] = i_icb_cmd_id ;
    end
    if(SPLT_PTR_1HOT == 1) begin:gen_ptr_1hot_rsp
        for(i = 0; i < SPLT_NUM; i = i+1)
        begin:gen_o_icb_rsp_ready
          assign o_icb_rsp_ready[i] = (o_icb_rsp_port_id[i] & i_icb_rsp_ready_pre);
        end
        assign i_icb_rsp_valid_pre = |(o_icb_rsp_valid & o_icb_rsp_port_id);
        reg sel_i_icb_rsp_err;
        reg sel_i_icb_rsp_excl_ok;
        reg [DW-1:0] sel_i_icb_rsp_rdata;
        reg [RSP_UW-1:0] sel_i_icb_rsp_usr;
        reg [ID_W-1:0] sel_i_icb_rsp_id;
        reg            sel_i_icb_rsp_last;
        always @ (*) begin : sel_icb_rsp_PROC
          sel_i_icb_rsp_err   = 1'b0;
          sel_i_icb_rsp_excl_ok   = 1'b0;
          sel_i_icb_rsp_rdata = {DW   {1'b0}};
          sel_i_icb_rsp_usr   = {RSP_UW{1'b0}};
          sel_i_icb_rsp_id   = {ID_W{1'b0}};
          sel_i_icb_rsp_last   = 1'b0;
          for(j = 0; j < SPLT_NUM; j = j+1) begin
            sel_i_icb_rsp_err     = sel_i_icb_rsp_err     | (       o_icb_rsp_port_id[j]   & o_icb_rsp_err[j]);
            sel_i_icb_rsp_excl_ok = sel_i_icb_rsp_excl_ok | (       o_icb_rsp_port_id[j]   & o_icb_rsp_excl_ok[j]);
            sel_i_icb_rsp_rdata   = sel_i_icb_rsp_rdata   | ({DW   {o_icb_rsp_port_id[j]}} & o_icb_rsp_rdata[j]);
            sel_i_icb_rsp_usr     = sel_i_icb_rsp_usr     | ({RSP_UW{o_icb_rsp_port_id[j]}} & o_icb_rsp_usr[j]);
            sel_i_icb_rsp_id      = sel_i_icb_rsp_id      | ({ID_W{o_icb_rsp_port_id[j]}} & o_icb_rsp_id[j]);
            sel_i_icb_rsp_last      = sel_i_icb_rsp_last      | (o_icb_rsp_port_id[j] & o_icb_rsp_last[j]);
          end
        end
        assign i_icb_rsp_err   = sel_i_icb_rsp_err  ;
        assign i_icb_rsp_excl_ok   = sel_i_icb_rsp_excl_ok  ;
        assign i_icb_rsp_rdata = sel_i_icb_rsp_rdata;
        assign i_icb_rsp_usr   = sel_i_icb_rsp_usr  ;
        assign i_icb_rsp_id    = sel_i_icb_rsp_id  ;
        assign i_icb_rsp_last    = sel_i_icb_rsp_last  ;
    end
    else begin:gen_ptr_not_1hot_rsp
        for(i = 0; i < SPLT_NUM; i = i+1)
        begin:gen_o_icb_rsp_ready
          assign o_icb_rsp_ready[i] = (o_icb_rsp_port_id == i[SPLT_PTR_W-1:0]) & i_icb_rsp_ready_pre;
        end
        assign i_icb_rsp_valid_pre = o_icb_rsp_valid[o_icb_rsp_port_id];
        assign i_icb_rsp_err     = o_icb_rsp_err    [o_icb_rsp_port_id];
        assign i_icb_rsp_excl_ok = o_icb_rsp_excl_ok[o_icb_rsp_port_id];
        assign i_icb_rsp_rdata   = o_icb_rsp_rdata  [o_icb_rsp_port_id];
        assign i_icb_rsp_usr     = o_icb_rsp_usr    [o_icb_rsp_port_id];
        assign i_icb_rsp_id     = o_icb_rsp_id    [o_icb_rsp_port_id];
        assign i_icb_rsp_last     = o_icb_rsp_last    [o_icb_rsp_port_id];
    end
  end
  endgenerate 
  assign splt_active = (i_icb_cmd_valid)
                     | (~rspid_fifo_empty)
                    ;
endmodule
module e603_subsys_gnrl_ficb_rw_splt_id # (
    parameter ID_W = 4,
  parameter ALLOW_DIFF = 1,
  parameter AW = 32,
  parameter DW = 32,
  parameter OUTS_FIFO_DP =4,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  input r_icb_support_oid,
  input w_icb_support_oid,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr,
  input                         icb_cmd_read,
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]              icb_cmd_wmask,
  input [CMD_UW-1:0]            icb_cmd_usr,
  input [ID_W-1:0]            icb_cmd_id,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [2:0]                   icb_cmd_size,
  input [7:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]           icb_rsp_usr,
  output [ID_W-1:0]           icb_rsp_id,
  output                      icb_rsp_last,
  input                         r_icb_cmd_ready,
  output                        r_icb_cmd_sel,
  output                        r_icb_cmd_valid,
  output[AW-1:0]                r_icb_cmd_addr,
  output                        r_icb_cmd_read,
  output[DW-1:0]                r_icb_cmd_wdata,
  output[DW/8-1:0]              r_icb_cmd_wmask,
  output[CMD_UW-1:0]            r_icb_cmd_usr,
  output[ID_W-1:0]            r_icb_cmd_id,
  output[1:0]                   r_icb_cmd_beat,
  output                        r_icb_cmd_lock,
  output                        r_icb_cmd_excl,
  output[2:0]                   r_icb_cmd_size,
  output[7:0]                   r_icb_cmd_xlen,
  output[1:0]                   r_icb_cmd_xburst,
  output[1:0]                   r_icb_cmd_modes,
  output                        r_icb_cmd_dmode,
  output[2:0]                   r_icb_cmd_attri,
  output                        r_icb_rsp_ready,
  input                         r_icb_rsp_valid,
  input                         r_icb_rsp_err  ,
  input                         r_icb_rsp_excl_ok,
  input  [DW-1:0]               r_icb_rsp_rdata,
  input  [RSP_UW-1:0]           r_icb_rsp_usr,
  input  [ID_W-1:0]           r_icb_rsp_id,
  input                       r_icb_rsp_last,
  input                         w_icb_cmd_ready,
  output                        w_icb_cmd_sel,
  output                        w_icb_cmd_valid,
  output[AW-1:0]                w_icb_cmd_addr,
  output                        w_icb_cmd_read,
  output[DW-1:0]                w_icb_cmd_wdata,
  output[DW/8-1:0]              w_icb_cmd_wmask,
  output[CMD_UW-1:0]            w_icb_cmd_usr,
  output[ID_W-1:0]            w_icb_cmd_id,
  output[1:0]                   w_icb_cmd_beat,
  output                        w_icb_cmd_lock,
  output                        w_icb_cmd_excl,
  output[2:0]                   w_icb_cmd_size,
  output[7:0]                   w_icb_cmd_xlen,
  output[1:0]                   w_icb_cmd_xburst,
  output[1:0]                   w_icb_cmd_modes,
  output                        w_icb_cmd_dmode,
  output[2:0]                   w_icb_cmd_attri,
  output                        w_icb_rsp_ready,
  input                         w_icb_rsp_valid,
  input                         w_icb_rsp_err  ,
  input                         w_icb_rsp_excl_ok,
  input  [DW-1:0]               w_icb_rsp_rdata,
  input  [RSP_UW-1:0]           w_icb_rsp_usr,
  input  [ID_W-1:0]           w_icb_rsp_id,
  input                       w_icb_rsp_last,
  input                         clk,
  input                         rst_n
  );
   wire [1:0] icb_cmd_splt_indic ={
      (~icb_cmd_read),
      icb_cmd_read
      };
  localparam SPLT_I_NUM = 2;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_sel;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_ready;
  wire [SPLT_I_NUM*AW-1:0] splt_bus_icb_cmd_addr;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_read;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_cmd_wdata;
  wire [SPLT_I_NUM*DW/8-1:0] splt_bus_icb_cmd_wmask;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_beat;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_lock;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_excl;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_size;
  wire [SPLT_I_NUM*CMD_UW-1:0] splt_bus_icb_cmd_usr;
  wire [SPLT_I_NUM*ID_W-1:0] splt_bus_icb_cmd_id;
  wire [SPLT_I_NUM*8-1:0] splt_bus_icb_cmd_xlen  ;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_xburst;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_modes ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_dmode ;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_attri ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_ready;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_err;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_excl_ok;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_rsp_rdata;
  wire [SPLT_I_NUM*RSP_UW-1:0] splt_bus_icb_rsp_usr;
  wire [SPLT_I_NUM*ID_W-1:0] splt_bus_icb_rsp_id;
  wire [SPLT_I_NUM-1:0] splt_bus_icb_rsp_last;
  assign {
                             w_icb_cmd_valid,
                             r_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
  assign {
                             w_icb_cmd_sel,
                             r_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
  assign {
                             w_icb_cmd_addr,
                             r_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
  assign {
                             w_icb_cmd_read,
                             r_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
  assign {
                             w_icb_cmd_wdata,
                             r_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
  assign {
                             w_icb_cmd_wmask,
                             r_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
  assign {
                             w_icb_cmd_xburst,
                             r_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
  assign {
                             w_icb_cmd_xlen,
                             r_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
  assign {
                             w_icb_cmd_modes,
                             r_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
  assign {
                             w_icb_cmd_dmode,
                             r_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
  assign {
                             w_icb_cmd_attri,
                             r_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
  assign {
                             w_icb_cmd_beat,
                             r_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
  assign {
                             w_icb_cmd_lock,
                             r_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
  assign {
                             w_icb_cmd_excl,
                             r_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
  assign {
                             w_icb_cmd_size,
                             r_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
  assign {
                             w_icb_cmd_usr,
                             r_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
  assign {
                             w_icb_cmd_id,
                             r_icb_cmd_id
                           } = splt_bus_icb_cmd_id;
  assign splt_bus_icb_cmd_ready = {
                             w_icb_cmd_ready,
                             r_icb_cmd_ready
                           };
  assign splt_bus_icb_rsp_valid = {
                             w_icb_rsp_valid,
                             r_icb_rsp_valid
                           };
  assign splt_bus_icb_rsp_err = {
                             w_icb_rsp_err,
                             r_icb_rsp_err
                           };
  assign splt_bus_icb_rsp_excl_ok = {
                             w_icb_rsp_excl_ok,
                             r_icb_rsp_excl_ok
                           };
  assign splt_bus_icb_rsp_rdata = {
                             w_icb_rsp_rdata,
                             r_icb_rsp_rdata
                           };
  assign splt_bus_icb_rsp_id = {
                             w_icb_rsp_id,
                             r_icb_rsp_id
                           };
  assign splt_bus_icb_rsp_last = {
                             w_icb_rsp_last,
                             r_icb_rsp_last
                           };
  assign splt_bus_icb_rsp_usr = {
                             w_icb_rsp_usr,
                             r_icb_rsp_usr
                           };
  assign {
                             w_icb_rsp_ready,
                             r_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
  e603_subsys_gnrl_ficb_splt_id # (
    .ID_W(ID_W),
  .USE_ALL_READY(0),
  .ALLOW_DIFF (ALLOW_DIFF),
  .ALLOW_0CYCL_RSP (0),
  .FIFO_OUTS_NUM   (OUTS_FIFO_DP),
  .FIFO_CUT_READY  (1),
  .SPLT_NUM   (2),
  .SPLT_PTR_W (2),
  .SPLT_PTR_1HOT (1),
  .CMD_UW     (CMD_UW),
  .RSP_UW     (RSP_UW),
  .AW         (AW),
  .DW         (DW)
  ) u_icb_rw_splt(
  .clk_en(1'b1),
  .splt_active            (),
  .i_icb_splt_indic       (icb_cmd_splt_indic),
  .o_icb_support_oid({w_icb_support_oid,r_icb_support_oid}),
  .i_icb_cmd_sel          (icb_cmd_sel )     ,
  .i_icb_cmd_valid        (icb_cmd_valid )     ,
  .i_icb_cmd_ready        (icb_cmd_ready )     ,
  .i_icb_cmd_read         (icb_cmd_read )      ,
  .i_icb_cmd_addr         (icb_cmd_addr )      ,
  .i_icb_cmd_wdata        (icb_cmd_wdata )     ,
  .i_icb_cmd_wmask        (icb_cmd_wmask)      ,
  .i_icb_cmd_beat         (icb_cmd_beat )     ,
  .i_icb_cmd_excl         (icb_cmd_excl )     ,
  .i_icb_cmd_lock         (icb_cmd_lock )     ,
  .i_icb_cmd_size         (icb_cmd_size )     ,
  .i_icb_cmd_xburst       (icb_cmd_xburst),
  .i_icb_cmd_xlen         (icb_cmd_xlen  ),
  .i_icb_cmd_modes        (icb_cmd_modes ),
  .i_icb_cmd_dmode        (icb_cmd_dmode ),
  .i_icb_cmd_attri        (icb_cmd_attri ),
  .i_icb_cmd_usr          (icb_cmd_usr   ),
  .i_icb_cmd_id          (icb_cmd_id   ),
  .i_icb_rsp_valid        (icb_rsp_valid )     ,
  .i_icb_rsp_ready        (icb_rsp_ready )     ,
  .i_icb_rsp_err          (icb_rsp_err)        ,
  .i_icb_rsp_excl_ok      (icb_rsp_excl_ok)    ,
  .i_icb_rsp_rdata        (icb_rsp_rdata )     ,
  .i_icb_rsp_usr          (icb_rsp_usr )     ,
  .i_icb_rsp_id          (icb_rsp_id )     ,
  .i_icb_rsp_last          (icb_rsp_last )     ,
  .o_bus_icb_cmd_ready    (splt_bus_icb_cmd_ready ) ,
  .o_bus_icb_cmd_valid    (splt_bus_icb_cmd_valid ) ,
  .o_bus_icb_cmd_sel      (splt_bus_icb_cmd_sel   ) ,
  .o_bus_icb_cmd_read     (splt_bus_icb_cmd_read )  ,
  .o_bus_icb_cmd_addr     (splt_bus_icb_cmd_addr )  ,
  .o_bus_icb_cmd_wdata    (splt_bus_icb_cmd_wdata ) ,
  .o_bus_icb_cmd_wmask    (splt_bus_icb_cmd_wmask)  ,
  .o_bus_icb_cmd_beat     (splt_bus_icb_cmd_beat ),
  .o_bus_icb_cmd_excl     (splt_bus_icb_cmd_excl ),
  .o_bus_icb_cmd_lock     (splt_bus_icb_cmd_lock ),
  .o_bus_icb_cmd_size     (splt_bus_icb_cmd_size ),
  .o_bus_icb_cmd_usr      (splt_bus_icb_cmd_usr  ),
  .o_bus_icb_cmd_id      (splt_bus_icb_cmd_id  ),
  .o_bus_icb_cmd_xburst   (splt_bus_icb_cmd_xburst),
  .o_bus_icb_cmd_xlen     (splt_bus_icb_cmd_xlen  ),
  .o_bus_icb_cmd_modes    (splt_bus_icb_cmd_modes ),
  .o_bus_icb_cmd_dmode    (splt_bus_icb_cmd_dmode ),
  .o_bus_icb_cmd_attri    (splt_bus_icb_cmd_attri ),
  .o_bus_icb_rsp_valid    (splt_bus_icb_rsp_valid ) ,
  .o_bus_icb_rsp_ready    (splt_bus_icb_rsp_ready ) ,
  .o_bus_icb_rsp_err      (splt_bus_icb_rsp_err)    ,
  .o_bus_icb_rsp_excl_ok  (splt_bus_icb_rsp_excl_ok),
  .o_bus_icb_rsp_rdata    (splt_bus_icb_rsp_rdata ) ,
  .o_bus_icb_rsp_usr      (splt_bus_icb_rsp_usr ) ,
  .o_bus_icb_rsp_id      (splt_bus_icb_rsp_id ) ,
  .o_bus_icb_rsp_last      (splt_bus_icb_rsp_last ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
`include "global.v"
module e603_subsys_gnrl_ficb_pd # (
  parameter AW = 32,
  parameter DW = 32,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter ASYNC_FF_LEVELS = 2,
  parameter OUTS_FIFO_DP =4,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1 
) (
  input              clk_en,
  input              i_icb_pd_n,
  input              i_icb_cmd_sel, 
  input              i_icb_cmd_valid, 
  output             i_icb_cmd_ready, 
  input              i_icb_cmd_read, 
  input  [AW-1:0]    i_icb_cmd_addr, 
  input  [DW-1:0]    i_icb_cmd_wdata, 
  input  [DW/8-1:0]  i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  output             i_icb_rsp_valid, 
  input              i_icb_rsp_ready, 
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [DW-1:0]    i_icb_rsp_rdata, 
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output             o_icb_cmd_sel, 
  output             o_icb_cmd_valid, 
  input              o_icb_cmd_ready, 
  output             o_icb_cmd_read, 
  output [AW-1:0]    o_icb_cmd_addr, 
  output [DW-1:0]    o_icb_cmd_wdata, 
  output [DW/8-1:0]  o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid, 
  output             o_icb_rsp_ready, 
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata, 
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  clk_aon,  
  input  clk,  
  input  rst_n
  );
  wire                        err_icb_cmd_ready;
  wire                        err_icb_cmd_sel;
  wire                        err_icb_cmd_valid;
  wire[AW-1:0]                err_icb_cmd_addr; 
  wire                        err_icb_cmd_read; 
  wire[DW-1:0]                err_icb_cmd_wdata;
  wire[DW/8-1:0]              err_icb_cmd_wmask;
  wire[CMD_UW-1:0]            err_icb_cmd_usr;
  wire[1:0]                   err_icb_cmd_beat;
  wire                        err_icb_cmd_lock;
  wire                        err_icb_cmd_excl;
  wire[2:0]                   err_icb_cmd_size;
  wire[7:0]                   err_icb_cmd_xlen;
  wire[1:0]                   err_icb_cmd_xburst;
  wire[1:0]                   err_icb_cmd_modes;
  wire                        err_icb_cmd_dmode;
  wire[2:0]                   err_icb_cmd_attri;
  wire                        err_icb_rsp_ready;
  wire                        err_icb_rsp_valid;
  wire                        err_icb_rsp_err     = 1'b1;
  wire                        err_icb_rsp_excl_ok = 1'b0;
  wire [DW-1:0]               err_icb_rsp_rdata   = {DW{1'b0}};
  wire [RSP_UW-1:0]           err_icb_rsp_usr     = {RSP_UW{1'b0}};
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_err_rsp_gen_stage(
    .i_vld(err_icb_cmd_valid & clk_en), 
    .i_rdy(err_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(err_icb_rsp_valid), 
    .o_rdy(err_icb_rsp_ready & clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
  wire icb_pd_n_synced;
  e603_subsys_gnrl_sync # (
  .DP(ASYNC_FF_LEVELS),
  .DW(1)
  ) u_pd_sync(
      .din_a    (i_icb_pd_n),
      .dout     (icb_pd_n_synced),
      .clk      (clk_aon),
      .rst_n    (rst_n) 
  );
  wire icb_pd_synced = ~icb_pd_n_synced;
  wire icb_drop = icb_pd_synced
                ;
   wire [1:0] i_icb_cmd_splt_indic ={
      icb_drop,
      (~icb_drop) 
      };
  localparam SPLT_I_NUM = 2;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_sel;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_ready;
  wire [SPLT_I_NUM*AW-1:0] splt_bus_icb_cmd_addr;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_read;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_cmd_wdata;
  wire [SPLT_I_NUM*DW/8-1:0] splt_bus_icb_cmd_wmask;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_beat;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_lock;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_excl;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_size;
  wire [SPLT_I_NUM*CMD_UW-1:0] splt_bus_icb_cmd_usr;
  wire [SPLT_I_NUM*8-1:0] splt_bus_icb_cmd_xlen  ;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_xburst;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_modes ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_dmode ;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_attri ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_ready;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_err;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_excl_ok;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_rsp_rdata;
  wire [SPLT_I_NUM*RSP_UW-1:0] splt_bus_icb_rsp_usr; 
  assign {
                             err_icb_cmd_valid,
                             o_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
  assign {
                             err_icb_cmd_sel,
                             o_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
  assign {
                             err_icb_cmd_addr,
                             o_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
  assign {
                             err_icb_cmd_read,
                             o_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
  assign {
                             err_icb_cmd_wdata,
                             o_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
  assign {
                             err_icb_cmd_wmask,
                             o_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
  assign {
                             err_icb_cmd_xburst,
                             o_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
  assign {
                             err_icb_cmd_xlen,
                             o_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
  assign {
                             err_icb_cmd_modes,
                             o_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
  assign {
                             err_icb_cmd_dmode,
                             o_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
  assign {
                             err_icb_cmd_attri,
                             o_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
  assign {
                             err_icb_cmd_beat,
                             o_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
  assign {
                             err_icb_cmd_lock,
                             o_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
  assign {
                             err_icb_cmd_excl,
                             o_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
  assign {
                             err_icb_cmd_size,
                             o_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
  assign {
                             err_icb_cmd_usr,
                             o_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
  assign splt_bus_icb_cmd_ready = {
                             err_icb_cmd_ready,
                             o_icb_cmd_ready
                           };
  assign splt_bus_icb_rsp_valid = {
                             err_icb_rsp_valid,
                             o_icb_rsp_valid
                           };
  assign splt_bus_icb_rsp_err = {
                             err_icb_rsp_err,
                             o_icb_rsp_err
                           };
  assign splt_bus_icb_rsp_excl_ok = {
                             err_icb_rsp_excl_ok,
                             o_icb_rsp_excl_ok
                           };
  assign splt_bus_icb_rsp_rdata = {
                             err_icb_rsp_rdata,
                             o_icb_rsp_rdata
                           };
  assign splt_bus_icb_rsp_usr = {
                             err_icb_rsp_usr,
                             o_icb_rsp_usr
                           };
  assign {
                             err_icb_rsp_ready,
                             o_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
  e603_subsys_gnrl_ficb_splt # (
  .USE_ALL_READY   (0),
  .ALLOW_DIFF      (0),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (OUTS_FIFO_DP),
  .FIFO_CUT_READY  (1),
  .SPLT_NUM        (2),
  .SPLT_PTR_W      (2),
  .SPLT_PTR_1HOT   (1),
  .CMD_UW     (CMD_UW),
  .RSP_UW     (RSP_UW),
  .AW         (AW),
  .DW         (DW) 
  ) u_icb_pd_splt(
  .clk_en(clk_en),
  .splt_active            (),
  .i_icb_splt_indic       (i_icb_cmd_splt_indic),        
  .i_icb_cmd_sel          (i_icb_cmd_sel )     ,
  .i_icb_cmd_valid        (i_icb_cmd_valid )     ,
  .i_icb_cmd_ready        (i_icb_cmd_ready )     ,
  .i_icb_cmd_read         (i_icb_cmd_read )      ,
  .i_icb_cmd_addr         (i_icb_cmd_addr )      ,
  .i_icb_cmd_wdata        (i_icb_cmd_wdata )     ,
  .i_icb_cmd_wmask        (i_icb_cmd_wmask)      ,
  .i_icb_cmd_beat         (i_icb_cmd_beat )     ,
  .i_icb_cmd_excl         (i_icb_cmd_excl )     ,
  .i_icb_cmd_lock         (i_icb_cmd_lock )     ,
  .i_icb_cmd_size         (i_icb_cmd_size )     ,
  .i_icb_cmd_xburst       (i_icb_cmd_xburst),
  .i_icb_cmd_xlen         (i_icb_cmd_xlen  ),
  .i_icb_cmd_modes        (i_icb_cmd_modes ),
  .i_icb_cmd_dmode        (i_icb_cmd_dmode ),
  .i_icb_cmd_attri        (i_icb_cmd_attri ),
  .i_icb_cmd_usr          (i_icb_cmd_usr   ),
  .i_icb_rsp_valid        (i_icb_rsp_valid )     ,
  .i_icb_rsp_ready        (i_icb_rsp_ready )     ,
  .i_icb_rsp_err          (i_icb_rsp_err)        ,
  .i_icb_rsp_excl_ok      (i_icb_rsp_excl_ok)    ,
  .i_icb_rsp_rdata        (i_icb_rsp_rdata )     ,
  .i_icb_rsp_usr          (i_icb_rsp_usr )     ,
  .o_bus_icb_cmd_ready    (splt_bus_icb_cmd_ready ) ,
  .o_bus_icb_cmd_valid    (splt_bus_icb_cmd_valid ) ,
  .o_bus_icb_cmd_sel      (splt_bus_icb_cmd_sel   ) ,
  .o_bus_icb_cmd_read     (splt_bus_icb_cmd_read )  ,
  .o_bus_icb_cmd_addr     (splt_bus_icb_cmd_addr )  ,
  .o_bus_icb_cmd_wdata    (splt_bus_icb_cmd_wdata ) ,
  .o_bus_icb_cmd_wmask    (splt_bus_icb_cmd_wmask)  ,
  .o_bus_icb_cmd_beat     (splt_bus_icb_cmd_beat ),
  .o_bus_icb_cmd_excl     (splt_bus_icb_cmd_excl ),
  .o_bus_icb_cmd_lock     (splt_bus_icb_cmd_lock ),
  .o_bus_icb_cmd_size     (splt_bus_icb_cmd_size ),
  .o_bus_icb_cmd_usr      (splt_bus_icb_cmd_usr  ),
  .o_bus_icb_cmd_xburst   (splt_bus_icb_cmd_xburst),
  .o_bus_icb_cmd_xlen     (splt_bus_icb_cmd_xlen  ),
  .o_bus_icb_cmd_modes    (splt_bus_icb_cmd_modes ),
  .o_bus_icb_cmd_dmode    (splt_bus_icb_cmd_dmode ),
  .o_bus_icb_cmd_attri    (splt_bus_icb_cmd_attri ),
  .o_bus_icb_rsp_valid    (splt_bus_icb_rsp_valid ) ,
  .o_bus_icb_rsp_ready    (splt_bus_icb_rsp_ready ) ,
  .o_bus_icb_rsp_err      (splt_bus_icb_rsp_err)    ,
  .o_bus_icb_rsp_excl_ok  (splt_bus_icb_rsp_excl_ok),
  .o_bus_icb_rsp_rdata    (splt_bus_icb_rsp_rdata ) ,
  .o_bus_icb_rsp_usr      (splt_bus_icb_rsp_usr ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
`include "global.v"
module e603_subsys_gnrl_ficb_pd_id # (
  parameter ID_W = 32,
  parameter AW = 32,
  parameter DW = 32,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter ASYNC_FF_LEVELS = 2,
  parameter OUTS_FIFO_DP =4,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1 
) (
  input              clk_en,
  input              i_icb_pd_n,
  input              i_icb_cmd_sel, 
  input              i_icb_cmd_valid, 
  output             i_icb_cmd_ready, 
  input              i_icb_cmd_read, 
  input  [AW-1:0]    i_icb_cmd_addr, 
  input  [DW-1:0]    i_icb_cmd_wdata, 
  input  [DW/8-1:0]  i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [2:0]       i_icb_cmd_size,
  input  [1:0]       i_icb_cmd_beat,
  input  [CMD_UW-1:0] i_icb_cmd_usr,
  input  [7:0]       i_icb_cmd_xlen,
  input  [1:0]       i_icb_cmd_xburst,
  input  [1:0]       i_icb_cmd_modes,
  input              i_icb_cmd_dmode,
  input  [2:0]       i_icb_cmd_attri,
  input  [ID_W-1:0] i_icb_cmd_id,
  output             i_icb_rsp_valid, 
  input              i_icb_rsp_ready, 
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [DW-1:0]    i_icb_rsp_rdata, 
  output [RSP_UW-1:0] i_icb_rsp_usr,
  output [ID_W-1:0] i_icb_rsp_id,
  output            i_icb_rsp_last,
  output             o_icb_cmd_sel, 
  output             o_icb_cmd_valid, 
  input              o_icb_cmd_ready, 
  output             o_icb_cmd_read, 
  output [AW-1:0]    o_icb_cmd_addr, 
  output [DW-1:0]    o_icb_cmd_wdata, 
  output [DW/8-1:0]  o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [2:0]       o_icb_cmd_size,
  output [1:0]       o_icb_cmd_beat,
  output [CMD_UW-1:0] o_icb_cmd_usr,
  output [ID_W-1:0] o_icb_cmd_id,
  output [7:0]       o_icb_cmd_xlen,
  output [1:0]       o_icb_cmd_xburst,
  output [1:0]       o_icb_cmd_modes,
  output             o_icb_cmd_dmode,
  output [2:0]       o_icb_cmd_attri,
  input              o_icb_rsp_valid, 
  output             o_icb_rsp_ready, 
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata, 
  input  [RSP_UW-1:0] o_icb_rsp_usr,
  input  [ID_W-1:0] o_icb_rsp_id,
  input             o_icb_rsp_last,
  input  clk_aon,  
  input  clk,  
  input  rst_n
  );
  wire                        err_icb_cmd_ready;
  wire                        err_icb_cmd_sel;
  wire                        err_icb_cmd_valid;
  wire[AW-1:0]                err_icb_cmd_addr; 
  wire                        err_icb_cmd_read; 
  wire[DW-1:0]                err_icb_cmd_wdata;
  wire[DW/8-1:0]              err_icb_cmd_wmask;
  wire[CMD_UW-1:0]            err_icb_cmd_usr;
  wire[ID_W-1:0]            err_icb_cmd_id;
  wire[1:0]                   err_icb_cmd_beat;
  wire                        err_icb_cmd_lock;
  wire                        err_icb_cmd_excl;
  wire[2:0]                   err_icb_cmd_size;
  wire[7:0]                   err_icb_cmd_xlen;
  wire[1:0]                   err_icb_cmd_xburst;
  wire[1:0]                   err_icb_cmd_modes;
  wire                        err_icb_cmd_dmode;
  wire[2:0]                   err_icb_cmd_attri;
  wire                        err_icb_rsp_ready;
  wire                        err_icb_rsp_valid;
  wire                        err_icb_rsp_err     = 1'b1;
  wire                        err_icb_rsp_excl_ok = 1'b0;
  wire [DW-1:0]               err_icb_rsp_rdata   = {DW{1'b0}};
  wire [RSP_UW-1:0]           err_icb_rsp_usr     = {RSP_UW{1'b0}};
  wire [ID_W-1:0]           err_icb_rsp_id     = {ID_W{1'b0}};
  wire                      err_icb_rsp_last     = 1'b0;
  e603_subsys_gnrl_pipe_stage # (
    .CUT_READY(1),
    .DP (1),
    .DW (1)
  ) u_err_rsp_gen_stage(
    .i_vld(err_icb_cmd_valid & clk_en), 
    .i_rdy(err_icb_cmd_ready), 
    .i_dat(1'b0),
    .o_vld(err_icb_rsp_valid), 
    .o_rdy(err_icb_rsp_ready & clk_en), 
    .o_dat(),
    .clk  (clk  )                     ,
    .rst_n(rst_n)
  );
  wire icb_pd_n_synced;
  e603_subsys_gnrl_sync # (
  .DP(ASYNC_FF_LEVELS),
  .DW(1)
  ) u_pd_sync(
      .din_a    (i_icb_pd_n),
      .dout     (icb_pd_n_synced),
      .clk      (clk_aon),
      .rst_n    (rst_n) 
  );
  wire icb_pd_synced = ~icb_pd_n_synced;
  wire icb_drop = icb_pd_synced
                ;
   wire [1:0] i_icb_cmd_splt_indic ={
      icb_drop,
      (~icb_drop) 
      };
   wire [1:0] o_icb_support_oid ={
      1'b0,
      1'b1 
      };
  localparam SPLT_I_NUM = 2;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_sel;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_ready;
  wire [SPLT_I_NUM*AW-1:0] splt_bus_icb_cmd_addr;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_read;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_cmd_wdata;
  wire [SPLT_I_NUM*DW/8-1:0] splt_bus_icb_cmd_wmask;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_beat;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_lock;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_excl;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_size;
  wire [SPLT_I_NUM*CMD_UW-1:0] splt_bus_icb_cmd_usr;
  wire [SPLT_I_NUM*ID_W-1:0] splt_bus_icb_cmd_id;
  wire [SPLT_I_NUM*8-1:0] splt_bus_icb_cmd_xlen  ;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_xburst;
  wire [SPLT_I_NUM*2-1:0] splt_bus_icb_cmd_modes ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_cmd_dmode ;
  wire [SPLT_I_NUM*3-1:0] splt_bus_icb_cmd_attri ;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_valid;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_ready;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_err;
  wire [SPLT_I_NUM*1-1:0] splt_bus_icb_rsp_excl_ok;
  wire [SPLT_I_NUM*DW-1:0] splt_bus_icb_rsp_rdata;
  wire [SPLT_I_NUM*RSP_UW-1:0] splt_bus_icb_rsp_usr; 
  wire [SPLT_I_NUM*ID_W-1:0] splt_bus_icb_rsp_id; 
  wire [SPLT_I_NUM-1:0] splt_bus_icb_rsp_last; 
  assign {
                             err_icb_cmd_valid,
                             o_icb_cmd_valid
                           } = splt_bus_icb_cmd_valid;
  assign {
                             err_icb_cmd_sel,
                             o_icb_cmd_sel
                           } = splt_bus_icb_cmd_sel;
  assign {
                             err_icb_cmd_addr,
                             o_icb_cmd_addr
                           } = splt_bus_icb_cmd_addr;
  assign {
                             err_icb_cmd_read,
                             o_icb_cmd_read
                           } = splt_bus_icb_cmd_read;
  assign {
                             err_icb_cmd_wdata,
                             o_icb_cmd_wdata
                           } = splt_bus_icb_cmd_wdata;
  assign {
                             err_icb_cmd_wmask,
                             o_icb_cmd_wmask
                           } = splt_bus_icb_cmd_wmask;
  assign {
                             err_icb_cmd_xburst,
                             o_icb_cmd_xburst
                           } = splt_bus_icb_cmd_xburst;
  assign {
                             err_icb_cmd_xlen,
                             o_icb_cmd_xlen
                           } = splt_bus_icb_cmd_xlen;
  assign {
                             err_icb_cmd_modes,
                             o_icb_cmd_modes
                           } = splt_bus_icb_cmd_modes;
  assign {
                             err_icb_cmd_dmode,
                             o_icb_cmd_dmode
                           } = splt_bus_icb_cmd_dmode;
  assign {
                             err_icb_cmd_attri,
                             o_icb_cmd_attri
                           } = splt_bus_icb_cmd_attri;
  assign {
                             err_icb_cmd_beat,
                             o_icb_cmd_beat
                           } = splt_bus_icb_cmd_beat;
  assign {
                             err_icb_cmd_lock,
                             o_icb_cmd_lock
                           } = splt_bus_icb_cmd_lock;
  assign {
                             err_icb_cmd_excl,
                             o_icb_cmd_excl
                           } = splt_bus_icb_cmd_excl;
  assign {
                             err_icb_cmd_size,
                             o_icb_cmd_size
                           } = splt_bus_icb_cmd_size;
  assign {
                             err_icb_cmd_usr,
                             o_icb_cmd_usr
                           } = splt_bus_icb_cmd_usr;
  assign {
                             err_icb_cmd_id,
                             o_icb_cmd_id
                           } = splt_bus_icb_cmd_id;
  assign splt_bus_icb_cmd_ready = {
                             err_icb_cmd_ready,
                             o_icb_cmd_ready
                           };
  assign splt_bus_icb_rsp_valid = {
                             err_icb_rsp_valid,
                             o_icb_rsp_valid
                           };
  assign splt_bus_icb_rsp_err = {
                             err_icb_rsp_err,
                             o_icb_rsp_err
                           };
  assign splt_bus_icb_rsp_excl_ok = {
                             err_icb_rsp_excl_ok,
                             o_icb_rsp_excl_ok
                           };
  assign splt_bus_icb_rsp_rdata = {
                             err_icb_rsp_rdata,
                             o_icb_rsp_rdata
                           };
  assign splt_bus_icb_rsp_usr = {
                             err_icb_rsp_usr,
                             o_icb_rsp_usr
                           };
  assign splt_bus_icb_rsp_id = {
                             err_icb_rsp_id,
                             o_icb_rsp_id
                           };
  assign splt_bus_icb_rsp_last = {
                             err_icb_rsp_last,
                             o_icb_rsp_last
                           };
  assign {
                             err_icb_rsp_ready,
                             o_icb_rsp_ready
                           } = splt_bus_icb_rsp_ready;
  e603_subsys_gnrl_ficb_splt_id # (
  .ID_W     (ID_W),
  .USE_ALL_READY   (0),
  .ALLOW_DIFF      (0),
  .ALLOW_0CYCL_RSP (ALLOW_0CYCL_RSP),
  .FIFO_OUTS_NUM   (OUTS_FIFO_DP),
  .FIFO_CUT_READY  (1),
  .SPLT_NUM        (2),
  .SPLT_PTR_W      (2),
  .SPLT_PTR_1HOT   (1),
  .CMD_UW     (CMD_UW),
  .RSP_UW     (RSP_UW),
  .AW         (AW),
  .DW         (DW) 
  ) u_icb_pd_splt(
  .clk_en(clk_en),
  .splt_active            (),
  .i_icb_splt_indic       (i_icb_cmd_splt_indic),        
  .o_icb_support_oid(o_icb_support_oid),
  .i_icb_cmd_sel          (i_icb_cmd_sel )     ,
  .i_icb_cmd_valid        (i_icb_cmd_valid )     ,
  .i_icb_cmd_ready        (i_icb_cmd_ready )     ,
  .i_icb_cmd_read         (i_icb_cmd_read )      ,
  .i_icb_cmd_addr         (i_icb_cmd_addr )      ,
  .i_icb_cmd_wdata        (i_icb_cmd_wdata )     ,
  .i_icb_cmd_wmask        (i_icb_cmd_wmask)      ,
  .i_icb_cmd_beat         (i_icb_cmd_beat )     ,
  .i_icb_cmd_excl         (i_icb_cmd_excl )     ,
  .i_icb_cmd_lock         (i_icb_cmd_lock )     ,
  .i_icb_cmd_size         (i_icb_cmd_size )     ,
  .i_icb_cmd_xburst       (i_icb_cmd_xburst),
  .i_icb_cmd_xlen         (i_icb_cmd_xlen  ),
  .i_icb_cmd_modes        (i_icb_cmd_modes ),
  .i_icb_cmd_dmode        (i_icb_cmd_dmode ),
  .i_icb_cmd_attri        (i_icb_cmd_attri ),
  .i_icb_cmd_usr          (i_icb_cmd_usr   ),
  .i_icb_cmd_id           (i_icb_cmd_id    ),
  .i_icb_rsp_valid        (i_icb_rsp_valid )     ,
  .i_icb_rsp_ready        (i_icb_rsp_ready )     ,
  .i_icb_rsp_err          (i_icb_rsp_err)        ,
  .i_icb_rsp_excl_ok      (i_icb_rsp_excl_ok)    ,
  .i_icb_rsp_rdata        (i_icb_rsp_rdata )     ,
  .i_icb_rsp_usr          (i_icb_rsp_usr )     ,
  .i_icb_rsp_id           (i_icb_rsp_id  )     ,
  .i_icb_rsp_last           (i_icb_rsp_last  )     ,
  .o_bus_icb_cmd_ready    (splt_bus_icb_cmd_ready ) ,
  .o_bus_icb_cmd_valid    (splt_bus_icb_cmd_valid ) ,
  .o_bus_icb_cmd_sel      (splt_bus_icb_cmd_sel   ) ,
  .o_bus_icb_cmd_read     (splt_bus_icb_cmd_read )  ,
  .o_bus_icb_cmd_addr     (splt_bus_icb_cmd_addr )  ,
  .o_bus_icb_cmd_wdata    (splt_bus_icb_cmd_wdata ) ,
  .o_bus_icb_cmd_wmask    (splt_bus_icb_cmd_wmask)  ,
  .o_bus_icb_cmd_beat     (splt_bus_icb_cmd_beat ),
  .o_bus_icb_cmd_excl     (splt_bus_icb_cmd_excl ),
  .o_bus_icb_cmd_lock     (splt_bus_icb_cmd_lock ),
  .o_bus_icb_cmd_size     (splt_bus_icb_cmd_size ),
  .o_bus_icb_cmd_usr      (splt_bus_icb_cmd_usr  ),
  .o_bus_icb_cmd_id       (splt_bus_icb_cmd_id   ),
  .o_bus_icb_cmd_xburst   (splt_bus_icb_cmd_xburst),
  .o_bus_icb_cmd_xlen     (splt_bus_icb_cmd_xlen  ),
  .o_bus_icb_cmd_modes    (splt_bus_icb_cmd_modes ),
  .o_bus_icb_cmd_dmode    (splt_bus_icb_cmd_dmode ),
  .o_bus_icb_cmd_attri    (splt_bus_icb_cmd_attri ),
  .o_bus_icb_rsp_valid    (splt_bus_icb_rsp_valid ) ,
  .o_bus_icb_rsp_ready    (splt_bus_icb_rsp_ready ) ,
  .o_bus_icb_rsp_err      (splt_bus_icb_rsp_err)    ,
  .o_bus_icb_rsp_excl_ok  (splt_bus_icb_rsp_excl_ok),
  .o_bus_icb_rsp_rdata    (splt_bus_icb_rsp_rdata ) ,
  .o_bus_icb_rsp_usr      (splt_bus_icb_rsp_usr ) ,
  .o_bus_icb_rsp_id       (splt_bus_icb_rsp_id  ) ,
  .o_bus_icb_rsp_last       (splt_bus_icb_rsp_last  ) ,
  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );
endmodule
`include "global.v"
module e603_subsys_gnrl_ficb2axi_ar_id # (
  parameter ID_W = 4,
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_UW = 1 
) (
  output                        ar_pend_active,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input                         icb_cmd_read, 
  input [AW-1:0]                icb_cmd_addr, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input [ID_W-1:0]              icb_cmd_id,
  input                         axi_arready,
  output                        axi_arvalid,
  output [AW-1:0]               axi_araddr,
  output [AXLEN_W-1:0]                  axi_arlen,
  output [CMD_SIZE_W-1:0]                  axi_arsize,
  output [1:0]                  axi_arburst,
  output                        axi_arlock,
  output [3:0]                  axi_arcache,
  output [2:0]                  axi_arprot,
  output [CMD_UW-1:0]            axi_aruser,
  output [ID_W-1:0]            axi_arid,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_W = AW+AXLEN_W+CMD_SIZE_W+1+2+4+3+CMD_UW+ID_W 
                    ;
  wire              i_arvalid;
  wire [AW-1:0]     i_araddr;
  wire [AXLEN_W-1:0]        i_arlen;
  wire [CMD_SIZE_W-1:0]        i_arsize;
  wire [1:0]        i_arburst;
  wire              i_arlock;
  wire [3:0]        i_arcache;
  wire [2:0]        i_arprot;
  wire [CMD_UW-1:0]  i_aruser;
  wire [ID_W-1:0]  i_arid;
  wire [PACK_W-1:0] i_axi_pack;
  wire [PACK_W-1:0] o_axi_pack;
  wire i_axi_vld;
  wire i_axi_rdy;
  wire o_axi_vld;
  wire o_axi_rdy;
  wire axi_ar_ready;
  wire burst_flag_r;
  wire burst_flag_en;
  wire burst_flag_set;
  wire burst_flag_clr;
  assign burst_flag_en = burst_flag_set || burst_flag_clr;
  assign axi_ar_ready = axi_arready;
  assign burst_flag_set = icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[0] & icb_clk_en;
  assign burst_flag_clr = burst_flag_r && icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[1] & icb_clk_en;
e603_subsys_gnrl_dfflr #(1) burst_flag_dfflr (burst_flag_en, burst_flag_set, burst_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign ar_pend_active = burst_flag_r;
  assign icb_cmd_ready = i_axi_rdy | burst_flag_r;
  assign i_arvalid = icb_cmd_valid & (~burst_flag_r);
  assign i_araddr   = icb_cmd_addr;
  assign i_arlen     = icb_cmd_xlen[AXLEN_W-1:0];
  assign i_arburst   = ((icb_cmd_xlen == {AXLEN_W{1'b0}}) & (icb_cmd_xburst[1:0] == 2'b0)) ? 2'b01 : icb_cmd_xburst[1:0];
  assign i_arsize    = icb_cmd_size;
  assign i_arlock    = icb_cmd_excl; 
  wire icb_cmd_mmode  = (icb_cmd_modes == 2'd0);
  wire icb_cmd_smode  = (icb_cmd_modes == 2'd2);
  wire icb_cmd_ifu    = icb_cmd_attri[0];
  wire icb_cmd_device = icb_cmd_attri[1];
  wire icb_cmd_nc     = icb_cmd_attri[2];
  assign i_arcache   =  (icb_cmd_device & icb_cmd_nc) ? 4'b1011 : 
                        icb_cmd_device ? 4'b0000 :
                        icb_cmd_nc     ? 4'b0011 : 4'b1111;
  assign i_arprot[0] = icb_cmd_mmode;
  assign i_arprot[1] = 1'b0; 
  assign i_arprot[2] = icb_cmd_ifu;
  assign i_aruser    = icb_cmd_usr;
  assign i_arid    = icb_cmd_id;
  assign i_axi_pack = 
                      {
                        i_araddr,
                        i_arlen,
                        i_arsize,
                        i_arburst,
                        i_arlock,
                        i_arcache,
                        i_arprot,
                        i_arid,
                        i_aruser 
                      };
  assign {
           axi_araddr,
           axi_arlen,
           axi_arsize,
           axi_arburst,
           axi_arlock,
           axi_arcache,
           axi_arprot,
           axi_arid,
           axi_aruser 
         } = o_axi_pack;
  assign axi_arvalid = o_axi_vld;
  assign i_axi_vld = i_arvalid;
  assign o_axi_rdy = axi_ar_ready;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_W)
  ) u_axi_ar_fifo (
        .i_clk_en(icb_clk_en),
        .i_vld(i_axi_vld),
        .i_rdy(i_axi_rdy),
        .i_dat(i_axi_pack),
        .o_clk_en(axi_bus_clk_en),
        .o_vld(o_axi_vld),
        .o_rdy(o_axi_rdy),  
        .o_dat(o_axi_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb2axi_aw_id # (
  parameter ID_W = 4,
  parameter SUPPORT_AWID_OOO = 0,
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_UW = 1
) (
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [ID_W -1:0]             icb_cmd_id,
  input                         axi_awready,
  output                        axi_awvalid,
  output [AW-1:0]               axi_awaddr,
  output [AXLEN_W-1:0]                  axi_awlen,
  output [CMD_SIZE_W-1:0]                  axi_awsize,
  output [1:0]                  axi_awburst,
  output                        axi_awlock,
  output [3:0]                  axi_awcache,
  output [2:0]                  axi_awprot,
  output [CMD_UW-1:0]            axi_awuser, 
  output [ID_W-1:0]            axi_awid, 
  input                         axi_wready,
  output                        axi_wvalid,
  output [DW-1:0]               axi_wdata,
  output [DW/8-1:0]               axi_wstrb,
  output                        axi_wlast,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_A_W = AW+AXLEN_W+CMD_SIZE_W+1+2+4+3+CMD_UW+ID_W 
                           ;
  localparam PACK_D_W = DW+DW/8+1;
  wire axi_aw_ready;
  wire axi_w_ready;
  wire burst_flag_r;
  wire burst_flag_en;
  wire burst_flag_set;
  wire burst_flag_clr;
  wire [PACK_A_W-1:0] i_axi_a_pack;
  wire [PACK_A_W-1:0] o_axi_a_pack;
  wire [PACK_D_W-1:0] i_axi_d_pack;
  wire [PACK_D_W-1:0] o_axi_d_pack;
  wire i_axi_a_vld;
  wire i_axi_a_rdy;
  wire o_axi_a_vld;
  wire o_axi_a_rdy;
  wire i_axi_d_vld;
  wire i_axi_d_rdy;
  wire o_axi_d_vld;
  wire o_axi_d_rdy;
  wire                i_awready;
  wire                i_awvalid;
  wire [AW-1:0]       i_awaddr;
  wire [AXLEN_W-1:0]          i_awlen;
  wire [CMD_SIZE_W-1:0]          i_awsize;
  wire [1:0]          i_awburst;
  wire                i_awlock;
  wire [3:0]          i_awcache;
  wire [2:0]          i_awprot;
  wire [ID_W-1:0]     i_awid; 
  wire [CMD_UW-1:0]    i_awuser; 
  wire                i_wready;
  wire                i_wvalid;
  wire [DW-1:0]       i_wdata;
  wire [DW/8-1:0]       i_wstrb;
  wire                i_wlast;
  assign axi_aw_ready = axi_awready ;
  assign axi_w_ready  = axi_wready  ;
  assign i_axi_a_pack = 
                      {
                        i_awaddr,
                        i_awlen,
                        i_awsize,
                        i_awburst,
                        i_awlock,
                        i_awcache,
                        i_awprot,
                        i_awid,
                        i_awuser  
                      };
  assign i_axi_a_vld = i_awvalid;
  assign i_awready = i_axi_a_rdy; 
  assign {
          axi_awaddr,
          axi_awlen,
          axi_awsize,
          axi_awburst,
          axi_awlock,
          axi_awcache,
          axi_awprot,
          axi_awid,
          axi_awuser  
         } = o_axi_a_pack;
  assign axi_awvalid = o_axi_a_vld;
  assign o_axi_a_rdy = axi_aw_ready;
  assign i_axi_d_pack = 
                      {
                       i_wdata,
                       i_wstrb,
                       i_wlast
                      };
  assign i_axi_d_vld = i_wvalid;
  assign i_wready    = i_axi_d_rdy; 
  assign {
          axi_wdata,
          axi_wstrb,
          axi_wlast
         } = o_axi_d_pack;
  assign axi_wvalid  = o_axi_d_vld;
  assign o_axi_d_rdy = axi_w_ready;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_A_W)
  ) u_axi_aw_fifo (
        .i_clk_en(icb_clk_en),
        .i_vld(i_axi_a_vld),
        .i_rdy(i_axi_a_rdy),
        .i_dat(i_axi_a_pack),
        .o_clk_en(axi_bus_clk_en),
        .o_vld(o_axi_a_vld),
        .o_rdy(o_axi_a_rdy),  
        .o_dat(o_axi_a_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_D_W)
  ) u_axi_w_fifo (
        .i_clk_en(icb_clk_en),
        .i_vld(i_axi_d_vld),
        .i_rdy(i_axi_d_rdy),
        .i_dat(i_axi_d_pack),
        .o_clk_en(axi_bus_clk_en),
        .o_vld(o_axi_d_vld),
        .o_rdy(o_axi_d_rdy),  
        .o_dat(o_axi_d_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  assign burst_flag_en = burst_flag_set || burst_flag_clr;
  assign burst_flag_set = icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[0] & icb_clk_en
                        ;
  assign burst_flag_clr = burst_flag_r && icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[1] & icb_clk_en;
e603_subsys_gnrl_dfflr #(1) burst_flag_dfflr (burst_flag_en, burst_flag_set, burst_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_cmd_ready =   (i_awready || burst_flag_r) && (i_wready);
  assign i_awvalid = icb_cmd_valid && (!burst_flag_r) && i_wready;
  assign i_wvalid  = icb_cmd_valid && (i_awready || burst_flag_r);
  assign i_awaddr   = icb_cmd_addr;
  assign i_awlen     = icb_cmd_xlen[AXLEN_W-1:0];
  assign i_awburst   = ((icb_cmd_xlen == {AXLEN_W{1'b0}}) & (icb_cmd_xburst[1:0] == 2'b0)) ? 2'b01 : icb_cmd_xburst[1:0];
  assign i_awsize    = icb_cmd_size;
  assign i_awlock    = icb_cmd_excl; 
  wire icb_cmd_mmode  = (icb_cmd_modes == 2'd0);
  wire icb_cmd_smode  = (icb_cmd_modes == 2'd2);
  wire icb_cmd_ifu    = icb_cmd_attri[0];
  wire icb_cmd_device = icb_cmd_attri[1];
  wire icb_cmd_nc     = icb_cmd_attri[2];
  assign i_awcache   =  (icb_cmd_device & icb_cmd_nc) ? 4'b0111 : 
                        icb_cmd_device ? 4'b0000 :
                          icb_cmd_nc     ? 4'b0011 : 4'b1111;
  assign i_awprot[0] = icb_cmd_mmode;
  assign i_awprot[1] = 1'b0; 
  assign i_awprot[2] = 1'b0;
  assign i_awuser    = icb_cmd_usr;
  generate
    if(SUPPORT_AWID_OOO == 1) begin: awid_ooo_is1
  assign i_awid      = icb_cmd_id;
    end
    else begin: awid_ooo_is0
  assign i_awid      = {ID_W{1'b0}};
    end
  endgenerate
  assign i_wdata     = icb_cmd_wdata;
  assign i_wstrb     = icb_cmd_wmask;   
  assign i_wlast    = ((icb_cmd_beat == 2'b00) && !burst_flag_r) || icb_cmd_beat[1];
endmodule
module e603_subsys_gnrl_ficb2axi_r_id # (
  parameter ID_W = 4,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter REG_OUT = 0,
  parameter RSP_UW = 1 
) (
  input                          icb_cmd_cnt_is_0,
  output                         icb_rrsp_valid,
  input                          icb_rrsp_ready,
  output [DW-1:0]                icb_rrsp_rdata,
  output                         icb_rrsp_err,
  output                         icb_rrsp_excl_ok,
  output [RSP_UW-1:0]            icb_rrsp_usr,
  output [ID_W -1:0]             icb_rrsp_id,
  output                         icb_rrsp_last,
  output                         axi_rready,
  input                          axi_rvalid,
  input [RSP_UW-1:0]              axi_ruser,
  input [DW-1:0]                 axi_rdata,
  input [1:0]                    axi_rresp,
  input                          axi_rlast,
  input [ID_W-1:0]               axi_rid,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_W = DW+2+1+RSP_UW+ID_W;
  wire                          o_rvalid;
  wire [DW-1:0]                 o_rdata;
  wire [RSP_UW-1:0]              o_rusr;
  wire [ID_W -1:0]              o_rid;
  wire [1:0]                    o_rresp;
  wire                          o_rlast;
  wire [PACK_W-1:0] i_axi_pack;
  wire [PACK_W-1:0] o_axi_pack;
  wire i_axi_vld;
  wire i_axi_rdy;
  wire o_axi_vld;
  wire o_axi_rdy;
  assign i_axi_pack = 
                      {
                        axi_rid,
                        axi_ruser,
                        axi_rdata,
                        axi_rresp,
                        axi_rlast 
                      };
  assign {
          o_rid,
          o_rusr,
          o_rdata,
          o_rresp,
          o_rlast 
         } = o_axi_pack;
  assign o_rvalid = o_axi_vld;
  assign icb_rrsp_valid = (~icb_cmd_cnt_is_0) & o_rvalid      ;
  assign o_axi_rdy      = (~icb_cmd_cnt_is_0) & icb_rrsp_ready;
  assign i_axi_vld = axi_rvalid ;
  assign axi_rready = i_axi_rdy;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .REG_OUT (REG_OUT),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_W)
  ) u_axi_r_fifo (
        .i_clk_en(axi_bus_clk_en),
        .i_vld(i_axi_vld),
        .i_rdy(i_axi_rdy),
        .i_dat(i_axi_pack),
        .o_clk_en(icb_clk_en),
        .o_vld(o_axi_vld),
        .o_rdy(o_axi_rdy),  
        .o_dat(o_axi_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  wire icb_rrsp_err_tmp     = o_rresp[1]   
                 ;
  assign icb_rrsp_err = icb_rrsp_err_tmp;
  wire icb_rrsp_excl_ok_tmp = (o_rresp == 2'b01);
  assign icb_rrsp_excl_ok = icb_rrsp_excl_ok_tmp;
  assign icb_rrsp_rdata   = o_rdata;
  assign icb_rrsp_usr     = o_rusr;
  assign icb_rrsp_id     = o_rid;
  assign icb_rrsp_last     = o_rlast;
endmodule
module e603_subsys_gnrl_ficb2axi_b_id # (
  parameter ID_W = 4,
  parameter SUPPORT_AWID_OOO = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter RSP_UW = 1,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2 
) (
  input                          wrsp_burst_fifo_o_vld,
  output                         icb_wrsp_valid,
  input                          icb_wrsp_ready,
  output                         icb_wrsp_err,
  output                         icb_wrsp_excl_ok,
  output [RSP_UW-1:0]             icb_wrsp_usr,
  output [ID_W-1:0]             icb_wrsp_id,
  output                        icb_wrsp_last,
  output                         axi_bready,
  input                          axi_bvalid,
  input [1:0]                    axi_bresp,
  input [RSP_UW-1:0]              axi_buser,
  input [ID_W-1:0]              axi_bid,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input [7:0]                   wrsp_xlen,
  output                        wrsp_last,
  input [ID_W-1:0] wrsp_id,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_W = 2+RSP_UW+ID_W;
  wire [ID_W-1:0]              o_bid;
  wire [RSP_UW-1:0]              o_busr;
  wire [1:0]                    o_bresp;
  wire o_burst = (wrsp_xlen != 8'b0);
  wire [PACK_W-1:0] i_axi_pack;
  wire [PACK_W-1:0] o_axi_pack;
  wire i_axi_vld;
  wire i_axi_rdy;
  wire o_axi_vld;
  wire o_axi_rdy;
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_r_nxt;
  wire       burst_cnt_ena;
  assign i_axi_pack = 
                      {
                        axi_bresp,
                        axi_bid, 
                        axi_buser 
                      };
  assign {
          o_bresp,
          o_bid, 
          o_busr 
         } = o_axi_pack;
  assign i_axi_vld = axi_bvalid ;
  assign axi_bready = i_axi_rdy;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_W)
  ) u_axi_b_fifo (
        .i_clk_en(axi_bus_clk_en),
        .i_vld(i_axi_vld),
        .i_rdy(i_axi_rdy),
        .i_dat(i_axi_pack),
        .o_clk_en(icb_clk_en),
        .o_vld(o_axi_vld),
        .o_rdy(o_axi_rdy),  
        .o_dat(o_axi_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  wire burst_first = (burst_cnt_r == 8'd0);
  assign burst_cnt_r_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_cnt_ena = o_burst && icb_wrsp_valid && icb_wrsp_ready & icb_clk_en;
  assign burst_last = (burst_cnt_r == wrsp_xlen) & (~burst_first);
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_r_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_wrsp_valid   = wrsp_last ? o_axi_vld : wrsp_burst_fifo_o_vld;
  assign o_axi_rdy = icb_wrsp_ready && wrsp_last;
  wire icb_wrsp_err_tmp     = wrsp_last ? (o_bresp[1] 
                                        ): 1'b0;
  assign icb_wrsp_err     = icb_wrsp_err_tmp;
  wire icb_wrsp_excl_ok_tmp = wrsp_last ? (o_bresp == 2'b01) : 1'b0;
  assign icb_wrsp_excl_ok = icb_wrsp_excl_ok_tmp;
  assign icb_wrsp_usr     = wrsp_last ? o_busr : {RSP_UW{1'b0}};
  generate
    if(SUPPORT_AWID_OOO == 1) begin: wrsp_id_ooo_is1
  assign icb_wrsp_id     = o_bid;
    end
    else begin: wrsp_id_ooo_is0
  assign icb_wrsp_id     = wrsp_id;
    end
  endgenerate
  assign icb_wrsp_last     = wrsp_last;
  assign wrsp_last = burst_last | (wrsp_xlen == 8'd0);
   endmodule
module e603_subsys_gnrl_ficb2axi_read_id # (
  parameter ID_W = 4,
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter REG_OUT = 0,
  parameter OUTS_CNT_W = 4,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  output icb2axi_read_pend_active,
  input                         axi_arready,
  output                        axi_arvalid,
  output [AW-1:0]               axi_araddr,
  output [AXLEN_W-1:0]                  axi_arlen,
  output [CMD_SIZE_W-1:0]                  axi_arsize,
  output [1:0]                  axi_arburst,
  output                        axi_arlock,
  output [3:0]                  axi_arcache,
  output [2:0]                  axi_arprot,
  output [CMD_UW-1:0]            axi_aruser,
  output [ID_W-1:0]            axi_arid,
  output                        axi_rready,
  input                         axi_rvalid,
  input [DW-1:0]                axi_rdata,
  input [RSP_UW-1:0]             axi_ruser,
  input [ID_W-1:0]             axi_rid,
  input [1:0]                   axi_rresp,
  input                         axi_rlast,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input [ID_W-1:0]             icb_cmd_id,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]            icb_rsp_usr,
  output [ID_W-1:0]            icb_rsp_id,
  output                       icb_rsp_last,
  input                         clk,
  input                         rst_n
  );
  localparam CNT_W = 8;
  wire outs_cnt_inc = icb_cmd_valid & icb_cmd_ready & icb_clk_en;
  wire outs_cnt_dec = icb_rsp_valid & icb_rsp_ready & icb_clk_en;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [CNT_W-1:0] outs_cnt_r;
  wire [CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_cmd_cnt_full = (outs_cnt_r == {CNT_W{1'b1}});
  wire icb_cmd_cnt_is_0 = (outs_cnt_r == {CNT_W{1'b0}});
  wire icb_cmd_valid_raw;
  wire icb_cmd_ready_raw;
  assign icb_cmd_valid_raw = (~icb_cmd_cnt_full) & icb_cmd_valid;
  assign icb_cmd_ready     = (~icb_cmd_cnt_full) & icb_cmd_ready_raw;
  wire ar_pend_active;
  assign icb2axi_read_pend_active = (~icb_cmd_cnt_is_0) | ar_pend_active | axi_arvalid;
 e603_subsys_gnrl_ficb2axi_ar_id # (
            .ID_W (ID_W),
            .AXLEN_W (AXLEN_W),
            .AW (AW),
            .DW (DW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP),
            .CMD_SIZE_W(CMD_SIZE_W),
            .CMD_UW (CMD_UW)
   ) u_icb2axi_ar(
            .ar_pend_active(ar_pend_active),
            .icb_cmd_valid (icb_cmd_valid_raw),
            .icb_cmd_ready (icb_cmd_ready_raw),
            .icb_cmd_addr (icb_cmd_addr), 
            .icb_cmd_sel  (icb_cmd_sel), 
            .icb_cmd_xlen(icb_cmd_xlen),
            .icb_cmd_xburst(icb_cmd_xburst),
            .icb_cmd_modes (icb_cmd_modes ),
            .icb_cmd_dmode (icb_cmd_dmode ),
            .icb_cmd_attri (icb_cmd_attri ),
            .icb_cmd_read (icb_cmd_read), 
            .icb_cmd_wdata (icb_cmd_wdata),
            .icb_cmd_wmask (icb_cmd_wmask),
            .icb_cmd_beat (icb_cmd_beat),
            .icb_cmd_lock (icb_cmd_lock),
            .icb_cmd_excl (icb_cmd_excl),
            .icb_cmd_size (icb_cmd_size),
            .icb_cmd_usr (icb_cmd_usr),
            .icb_cmd_id  (icb_cmd_id ),
            .axi_arready (axi_arready),
            .axi_arvalid (axi_arvalid),
            .axi_araddr (axi_araddr),
            .axi_arlen (axi_arlen),
            .axi_arsize (axi_arsize),
            .axi_arburst (axi_arburst),
            .axi_arlock (axi_arlock),
            .axi_arcache (axi_arcache),
            .axi_arprot (axi_arprot),
            .axi_aruser (axi_aruser),
            .axi_arid (axi_arid),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .clk (clk),
            .rst_n (rst_n)
  );
  e603_subsys_gnrl_ficb2axi_r_id # (
            .ID_W (ID_W),
            .AW (AW),
            .DW (DW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP),
            .REG_OUT(REG_OUT),
            .RSP_UW (RSP_UW) 
  ) u_icb2axi_r(
            .icb_cmd_cnt_is_0(icb_cmd_cnt_is_0),
            .icb_rrsp_valid (icb_rsp_valid),
            .icb_rrsp_ready (icb_rsp_ready),
            .icb_rrsp_rdata (icb_rsp_rdata),
            .icb_rrsp_usr (icb_rsp_usr),
            .icb_rrsp_id (icb_rsp_id),
            .icb_rrsp_last (icb_rsp_last),
            .icb_rrsp_err (icb_rsp_err),
            .icb_rrsp_excl_ok (icb_rsp_excl_ok),
            .axi_rready (axi_rready),
            .axi_rvalid (axi_rvalid),
            .axi_rdata (axi_rdata),
            .axi_ruser (axi_ruser),
            .axi_rid (axi_rid),
            .axi_rresp (axi_rresp),
            .axi_rlast (axi_rlast),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .clk (clk),
            .rst_n (rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb2axi_write_id # (
  parameter ID_W = 4,
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter OUTS_CNT_W =2,
  parameter SUPPORT_AWID_OOO = 0,
  parameter OUTS_FIFO_DP =4,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP =2,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  output                        icb2axi_write_pend_active,
  input                         axi_awready,
  output                        axi_awvalid,
  output [AW-1:0]               axi_awaddr,
  output [AXLEN_W-1:0]                  axi_awlen,
  output [CMD_SIZE_W-1:0]                  axi_awsize,
  output [1:0]                  axi_awburst,
  output                        axi_awlock,
  output [3:0]                  axi_awcache,
  output [2:0]                  axi_awprot,
  output [CMD_UW-1:0]            axi_awuser, 
  output [ID_W-1:0]            axi_awid, 
  input                         axi_wready,
  output                        axi_wvalid,
  output [DW-1:0]               axi_wdata,
  output [DW/8-1:0]               axi_wstrb,
  output                        axi_wlast,
  output                         axi_bready,
  input                          axi_bvalid,
  input [RSP_UW-1:0]              axi_buser,
  input [ID_W-1:0]              axi_bid,
  input [1:0]                    axi_bresp,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr,
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input [ID_W-1:0]              icb_cmd_id,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err,
  output                        icb_rsp_excl_ok,
  output[RSP_UW-1:0]             icb_rsp_usr,
  output[DW-1:0]                icb_rsp_rdata,
  output[ID_W-1:0]              icb_rsp_id,
  output                        icb_rsp_last,
  input                         clk,
  input                         rst_n
  );
  assign icb_rsp_rdata = {DW{1'b0}};
  wire [7:0] wrsp_xlen;
  wire [7:0] wcmd_xlen;
  wire wrsp_burst_fifo_i_vld;
  wire wrsp_burst_fifo_o_rdy;
  wire wrsp_burst_fifo_o_vld;
  wire wrsp_burst_fifo_i_rdy;
  wire wrsp_last;
  wire icb_cmd_valid_raw;
  wire icb_cmd_ready_raw;
  assign icb_cmd_valid_raw = wrsp_burst_fifo_i_rdy & icb_cmd_valid;
  assign icb_cmd_ready     = wrsp_burst_fifo_i_rdy & icb_cmd_ready_raw;
  assign wrsp_burst_fifo_i_vld = icb_cmd_valid & icb_cmd_ready;
  assign wrsp_burst_fifo_o_rdy = icb_rsp_valid & icb_rsp_ready;
  assign wcmd_xlen = icb_cmd_xlen[7:0];
  wire [ID_W-1:0] wrsp_id;
  generate
    if(SUPPORT_AWID_OOO == 1) begin: ooo_is1
  assign wrsp_id = {ID_W{1'b0}};
  e603_subsys_ficbficb2axi_gnrl_ooo_id_buf # (
        .DP  (OUTS_FIFO_DP),
        .IDW(ID_W),
        .DP_PTR_W(OUTS_CNT_W),
        .DW  (8)
  ) u_wrsp_burst_ooo_id_buf (
        .i_vld(wrsp_burst_fifo_i_vld & icb_clk_en),
        .i_rdy(wrsp_burst_fifo_i_rdy),
        .i_id(icb_cmd_id),
        .o_id(icb_rsp_id),
        .o_match(),
        .i_dat(wcmd_xlen),
        .o_vld(wrsp_burst_fifo_o_vld),
        .o_rdy(wrsp_burst_fifo_o_rdy & icb_clk_en),  
        .o_dat(wrsp_xlen),  
        .clk  (clk),
        .rst_n(rst_n)
  );
    end
    else begin: ooo_is0
     e603_subsys_gnrl_fifo # (
        .REG_OUT(1),
        .DP  (OUTS_FIFO_DP),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DW  (
               ID_W+8)
  ) u_wrsp_burst_fifo (
        .i_vld(wrsp_burst_fifo_i_vld & icb_clk_en),
        .i_rdy(wrsp_burst_fifo_i_rdy),
        .i_dat({
            icb_cmd_id, wcmd_xlen}),
        .o_vld(wrsp_burst_fifo_o_vld),
        .o_rdy(wrsp_burst_fifo_o_rdy & icb_clk_en),  
        .o_dat({
            wrsp_id, wrsp_xlen}),  
        .clk  (clk),
        .rst_n(rst_n)
  );
    end
  endgenerate
 e603_subsys_gnrl_ficb2axi_aw_id # (
            .ID_W (ID_W),
            .SUPPORT_AWID_OOO (SUPPORT_AWID_OOO),
            .AXLEN_W (AXLEN_W),
            .AW (AW),
            .DW (DW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP),
            .CMD_SIZE_W(CMD_SIZE_W),
            .CMD_UW (CMD_UW) 
) u_icb2axi_aw (
            .icb_cmd_valid (icb_cmd_valid_raw),
            .icb_cmd_ready (icb_cmd_ready_raw),
            .icb_cmd_addr (icb_cmd_addr), 
            .icb_cmd_xlen(icb_cmd_xlen),
            .icb_cmd_xburst(icb_cmd_xburst),
            .icb_cmd_modes (icb_cmd_modes ),
            .icb_cmd_dmode (icb_cmd_dmode ),
            .icb_cmd_attri (icb_cmd_attri ),
            .icb_cmd_read (icb_cmd_read), 
            .icb_cmd_wdata (icb_cmd_wdata),
            .icb_cmd_wmask (icb_cmd_wmask),
            .icb_cmd_beat (icb_cmd_beat),
            .icb_cmd_lock (icb_cmd_lock),
            .icb_cmd_excl (icb_cmd_excl),
            .icb_cmd_size (icb_cmd_size),
            .icb_cmd_usr (icb_cmd_usr),
            .icb_cmd_id (icb_cmd_id),
            .axi_awready (axi_awready),
            .axi_awvalid (axi_awvalid),
            .axi_awaddr (axi_awaddr),
            .axi_awlen (axi_awlen),
            .axi_awsize (axi_awsize),
            .axi_awburst (axi_awburst),
            .axi_awlock (axi_awlock),
            .axi_awcache (axi_awcache),
            .axi_awprot (axi_awprot),
            .axi_awuser (axi_awuser),
            .axi_awid (axi_awid),
            .axi_wready (axi_wready),
            .axi_wvalid (axi_wvalid),
            .axi_wdata (axi_wdata),
            .axi_wstrb (axi_wstrb),
            .axi_wlast (axi_wlast),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .clk (clk),
            .rst_n (rst_n)
  );
  e603_subsys_gnrl_ficb2axi_b_id # (
            .ID_W (ID_W),
            .SUPPORT_AWID_OOO (SUPPORT_AWID_OOO),
            .AW (AW),
            .DW (DW),
            .RSP_UW (RSP_UW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP) 
   ) u_icb2axi_b(
            .wrsp_burst_fifo_o_vld (wrsp_burst_fifo_o_vld),
            .icb_wrsp_valid (icb_rsp_valid),
            .icb_wrsp_ready (icb_rsp_ready),
            .icb_wrsp_err (icb_rsp_err),
            .icb_wrsp_excl_ok (icb_rsp_excl_ok),
            .icb_wrsp_usr (icb_rsp_usr),
            .icb_wrsp_id (icb_rsp_id),
            .icb_wrsp_last (icb_rsp_last),
            .axi_bready (axi_bready),
            .axi_bvalid (axi_bvalid),
            .axi_bresp (axi_bresp),
            .axi_buser (axi_buser),
            .axi_bid (axi_bid),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .wrsp_xlen  (wrsp_xlen),
            .wrsp_last  (wrsp_last),
            .wrsp_id    (wrsp_id  ),
            .clk (clk),
            .rst_n (rst_n)
  );
  assign icb2axi_write_pend_active = wrsp_burst_fifo_o_vld | axi_wvalid | axi_awvalid;
endmodule
`include "global.v"
module e603_subsys_ficbficb2axi_gnrl_ooo_id_buf # (
  parameter IDW   = 32,
  parameter DP   = 8,
  parameter DP_PTR_W = 4,
  parameter DW   = 32
) (
  input           i_vld, 
  output          i_rdy, 
  input [IDW-1:0] i_id, 
  input  [DW-1:0] i_dat,
  output          o_vld, 
  output          o_match, 
  input           o_rdy, 
  output [DW-1:0] o_dat,
  input [IDW-1:0] o_id,  
  input           clk,
  input           rst_n
);
genvar i;
integer j;
    wire [DW-1:0] fifo_rf_r [DP-1:0];
    wire [IDW-1:0] fifo_id_r  [DP-1:0];
    wire [DP-1:0]  fifo_vld_set;
    wire [DP-1:0]  fifo_vld_clr;
    wire [DP-1:0]  fifo_vld_ena;
    wire [DP-1:0]  fifo_vld_nxt;
    wire [DP-1:0]  fifo_vld_r;
    wire [DP-1:0]  fifo_dep_set;
    wire [DP-1:0]  fifo_dep_clr;
    wire [DP-1:0]  fifo_dep_ena;
    wire [DP-1:0]  fifo_dep_nxt;
    wire [DP-1:0]  fifo_dep_r;
    wire [DP-1:0]  fifo_last_set;
    wire [DP-1:0]  fifo_last_clr;
    wire [DP-1:0]  fifo_last_ena;
    wire [DP-1:0]  fifo_last_nxt;
    wire [DP-1:0]  fifo_last_r;
    wire [DP_PTR_W-1:0] fifo_dep_entid_r [DP-1:0];
    wire [DP-1:0] fifo_rf_ena;
    wire wen = i_vld & i_rdy;
    wire ren = o_vld & o_rdy;
    wire [DP-1:0] rptr_vec_r;
    wire [DP-1:0] wptr_vec_r;
    wire [DP-1:0] i_id_match_id;
    wire [DP-1:0] i_id_match_id_noclr;
    wire [DP-1:0] i_id_match_id_last;
    reg [DP_PTR_W-1:0] i_id_match_id_entid;
  generate 
    for (i=0; i<DP; i=i+1) begin:gen_wptr_vec
      if(i == 0) begin: i_is_0
          assign wptr_vec_r[i] = (~fifo_vld_r[i]);
      end
      else begin: i_is_not0
          assign wptr_vec_r[i] = (~fifo_vld_r[i]) & (&fifo_vld_r[i-1:0]);
      end
      assign rptr_vec_r[i] = (fifo_vld_r[i] & (o_id == fifo_id_r[i]) & (~fifo_dep_r[i]));
      assign i_id_match_id[i] = (fifo_vld_r[i] & (i_id == fifo_id_r[i]));
      assign i_id_match_id_noclr[i] = i_id_match_id[i] & (~fifo_vld_clr[i]) ;
      assign i_id_match_id_last[i]  = i_id_match_id[i] & fifo_last_r[i] ;
    end
  endgenerate
      assign i_rdy = |(~fifo_vld_r);
  generate 
    for (i=0; i<DP; i=i+1) begin:gen_fifo_rf
      assign fifo_rf_ena[i] = wen & wptr_vec_r[i];
e603_subsys_gnrl_dfflr  #(DW) fifo_rf_dffl (fifo_rf_ena[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(IDW) fifo_id_dffl (fifo_rf_ena[i], i_id , fifo_id_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      assign fifo_vld_set[i] = fifo_rf_ena[i];
      assign fifo_vld_clr[i] = ren & rptr_vec_r[i];
      assign fifo_vld_ena[i] = fifo_vld_set[i] | fifo_vld_clr[i] ;
      assign fifo_vld_nxt[i] = fifo_vld_set[i];
e603_subsys_gnrl_dfflr #(1)  fifo_vld_dfflr (fifo_vld_ena[i], fifo_vld_nxt[i], fifo_vld_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      assign fifo_dep_set[i] = fifo_vld_set[i] & 
                                  (|i_id_match_id_noclr);
// spyglass disable_block ImproperRangeIndex-ML
// SMD: Index fifo_dep_entid_r of width is larger than the width required for the max value of the signal fifo_vld_clr
// SJ:  This is not cared
      assign fifo_dep_clr[i] = fifo_vld_clr[i] | (fifo_dep_r[i] & fifo_vld_clr[fifo_dep_entid_r[i]]);
// spyglass enable_block ImproperRangeIndex-ML
      assign fifo_dep_ena[i] = fifo_dep_set[i] | fifo_dep_clr[i] ;
      assign fifo_dep_nxt[i] = fifo_dep_set[i];
e603_subsys_gnrl_dfflr #(1)  fifo_dep_dffl (fifo_dep_ena[i], fifo_dep_nxt[i], fifo_dep_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      assign fifo_last_set[i] = fifo_vld_set[i]; 
      assign fifo_last_clr[i] = fifo_vld_clr[i] | (fifo_last_r[i] & wen & i_id_match_id[i]);
      assign fifo_last_ena[i] = fifo_last_set[i] | fifo_last_clr[i] ;
      assign fifo_last_nxt[i] = fifo_last_set[i];
e603_subsys_gnrl_dfflr #(1)  fifo_last_dffl (fifo_last_ena[i], fifo_last_nxt[i], fifo_last_r[i], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(DP_PTR_W)              fifo_dep_entid_dffl (fifo_dep_set[i], i_id_match_id_entid, fifo_dep_entid_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
  endgenerate
    always @*
        begin : fifo_dep_entid_nxt_PROC
          i_id_match_id_entid = {DP_PTR_W{1'b0}};
          for(j=0; j<DP; j=j+1) begin
// spyglass disable_block W216
// SMD: Inappropriate range select for int_part_sel variable
// SJ:  Here is not a real issue
            i_id_match_id_entid = i_id_match_id_entid | ({DP_PTR_W{i_id_match_id_last[j]}} & j[DP_PTR_W-1:0]);
// spyglass enable_block W216
          end
        end
    wire [DW-1:0] mux_rdat;
    reg [DW-1:0] mux_rdat_t;
        always @*
        begin : rd_port_PROC
          mux_rdat_t = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_t = mux_rdat_t | ({DW{rptr_vec_r[j]}} & fifo_rf_r[j]);
          end
        end
    assign mux_rdat = mux_rdat_t;
        assign o_dat = mux_rdat;
    assign o_vld = |fifo_vld_r;
    assign o_match = |rptr_vec_r;
endmodule 
module e603_subsys_gnrl_ficb2axi_read_async_id # (
  parameter ID_W = 4,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter OUTS_CNT_W = 4,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 1,
  parameter ASYNC_FIFO_DP = 6,
  parameter ASYNC_FIFO_DP_PTR_W = 3,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  output                        icb2axi_read_async_icb_active,
  output                        icb2axi_read_async_axi_active,
  output                        icb2axi_read_pend_active,
  input                         axi_arready,
  output                        axi_arvalid,
  output [AW-1:0]               axi_araddr,
  output [7:0]                  axi_arlen,
  output [CMD_SIZE_W-1:0]                  axi_arsize,
  output [1:0]                  axi_arburst,
  output                        axi_arlock,
  output [3:0]                  axi_arcache,
  output [2:0]                  axi_arprot,
  output [CMD_UW-1:0]            axi_aruser,
  output [ID_W-1:0]            axi_arid,
  output                        axi_rready,
  input                         axi_rvalid,
  input [DW-1:0]                axi_rdata,
  input [RSP_UW-1:0]             axi_ruser,
  input [ID_W-1:0]             axi_rid,
  input [1:0]                   axi_rresp,
  input                         axi_rlast,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [7:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input [ID_W-1:0]             icb_cmd_id,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]            icb_rsp_usr,
  output [ID_W-1:0]            icb_rsp_id,
  output                       icb_rsp_last,
  input  async_axi_clk,
  input  async_axi_rst_n,
  input  icb_clk,
  input  icb_rst_n
  );
  wire i_icb_reset_flag_r;
e603_subsys_gnrl_dffrs #(1) reset_flag_dffrs (1'b0, i_icb_reset_flag_r, icb_clk, icb_rst_n);// VPP_NO_REG_PARSE
  wire i_icb_cmd_valid;
  wire i_icb_cmd_ready;
  assign i_icb_cmd_valid = (~i_icb_reset_flag_r) & icb_cmd_valid;
  assign icb_cmd_ready   = (~i_icb_reset_flag_r) & i_icb_cmd_ready;
  wire                        icb2axi_arready;
  wire                        icb2axi_arvalid;
  wire [AW-1:0]               icb2axi_araddr;
  wire [7:0]                  icb2axi_arlen;
  wire [CMD_SIZE_W-1:0]                  icb2axi_arsize;
  wire [1:0]                  icb2axi_arburst;
  wire                        icb2axi_arlock;
  wire [3:0]                  icb2axi_arcache;
  wire [2:0]                  icb2axi_arprot;
  wire [CMD_UW-1:0]           icb2axi_aruser;
  wire [ID_W-1:0]           icb2axi_arid;
  localparam AR_PACK_W = (AW+8+CMD_SIZE_W+2+1+4+3+CMD_UW+ID_W) 
          ;
  wire [AR_PACK_W-1:0] ar_fifo_i_dat = {
                              icb2axi_araddr,
                              icb2axi_arlen,
                              icb2axi_arsize,
                              icb2axi_arburst,
                              icb2axi_arlock,
                              icb2axi_arcache,
                              icb2axi_arprot,
                              icb2axi_arid, 
                              icb2axi_aruser 
                                 };
  wire [AR_PACK_W-1:0] ar_fifo_o_dat;
  assign {
                              axi_araddr,
                              axi_arlen,
                              axi_arsize,
                              axi_arburst,
                              axi_arlock,
                              axi_arcache,
                              axi_arprot,
                              axi_arid,
                              axi_aruser
                                } = ar_fifo_o_dat;
  wire                        icb2axi_rready;
  wire                        icb2axi_rvalid;
  wire[DW-1:0]                icb2axi_rdata;
  wire[RSP_UW-1:0]            icb2axi_ruser;
  wire[ID_W-1:0]              icb2axi_rid;
  wire[1:0]                   icb2axi_rresp;
  wire                        icb2axi_rlast;
  localparam R_PACK_W = (1+2+DW+RSP_UW+ID_W);
  wire [R_PACK_W-1:0] r_fifo_i_dat = {
                              axi_rdata,
                              axi_ruser,
                              axi_rid,
                              axi_rresp,
                              axi_rlast 
                                 };
  wire [R_PACK_W-1:0] r_fifo_o_dat;
  assign {
                              icb2axi_rdata,
                              icb2axi_ruser,
                              icb2axi_rid,
                              icb2axi_rresp,
                              icb2axi_rlast 
                                 } = r_fifo_o_dat;
wire i_icb2axi_read_pend_active;
 e603_subsys_gnrl_ficb2axi_read_id # (
            .ID_W (ID_W),
            .AW (AW),
            .DW (DW),
            .OUTS_CNT_W(OUTS_CNT_W),
            .RATIO_FIFO_DP(0),
            .CMD_UW (CMD_UW),
            .RSP_UW (RSP_UW)
   ) u_icb2axi_read(
            .icb2axi_read_pend_active(i_icb2axi_read_pend_active),
            .icb_cmd_valid    (i_icb_cmd_valid),
            .icb_cmd_ready    (i_icb_cmd_ready),
            .icb_cmd_addr     (icb_cmd_addr), 
            .icb_cmd_sel      (icb_cmd_sel), 
            .icb_cmd_xlen     (icb_cmd_xlen),
            .icb_cmd_xburst   (icb_cmd_xburst),
            .icb_cmd_modes    (icb_cmd_modes ),
            .icb_cmd_dmode    (icb_cmd_dmode ),
            .icb_cmd_attri    (icb_cmd_attri ),
            .icb_cmd_read     (icb_cmd_read), 
            .icb_cmd_wdata    (icb_cmd_wdata),
            .icb_cmd_wmask    (icb_cmd_wmask),
            .icb_cmd_beat     (icb_cmd_beat),
            .icb_cmd_lock     (icb_cmd_lock),
            .icb_cmd_excl     (icb_cmd_excl),
            .icb_cmd_size     (icb_cmd_size),
            .icb_cmd_usr      (icb_cmd_usr),
            .icb_cmd_id       (icb_cmd_id ),
            .icb_rsp_valid   (icb_rsp_valid),
            .icb_rsp_ready   (icb_rsp_ready),
            .icb_rsp_rdata   (icb_rsp_rdata),
            .icb_rsp_usr     (icb_rsp_usr),
            .icb_rsp_err     (icb_rsp_err),
            .icb_rsp_excl_ok (icb_rsp_excl_ok),
            .icb_rsp_id     (icb_rsp_id),
            .icb_rsp_last     (icb_rsp_last),
            .axi_arready (icb2axi_arready),
            .axi_arvalid (icb2axi_arvalid),
            .axi_araddr  (icb2axi_araddr),
            .axi_arlen   (icb2axi_arlen),
            .axi_arsize  (icb2axi_arsize),
            .axi_arburst (icb2axi_arburst),
            .axi_arlock  (icb2axi_arlock),
            .axi_arcache (icb2axi_arcache),
            .axi_arprot  (icb2axi_arprot),
            .axi_aruser  (icb2axi_aruser),
            .axi_arid  (icb2axi_arid),
            .axi_rready (icb2axi_rready),
            .axi_rvalid (icb2axi_rvalid),
            .axi_rdata  (icb2axi_rdata),
            .axi_ruser  (icb2axi_ruser),
            .axi_rid  (icb2axi_rid),
            .axi_rresp  (icb2axi_rresp),
            .axi_rlast  (icb2axi_rlast),
            .axi_bus_clk_en (1'b1),
            .icb_clk_en (1'b1),
            .clk   (icb_clk),
            .rst_n (icb_rst_n) 
  );
  wire ar_async_i_active;
  wire ar_async_o_active;
  wire r_async_i_active;
  wire r_async_o_active;
  e603_subsys_gnrl_cdc_fifo # (
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (AR_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_ar(
    .i_clk   (icb_clk),
    .i_rst_n (icb_rst_n),
    .o_clk   (async_axi_clk),
    .o_rst_n (async_axi_rst_n),
    .i_vld    (icb2axi_arvalid),
    .i_rdy    (icb2axi_arready),
    .i_dat    (ar_fifo_i_dat),
    .i_cdc_fifo_active(ar_async_i_active),
    .o_cdc_fifo_active(ar_async_o_active),
    .o_vld    (axi_arvalid),
    .o_rdy    (axi_arready),
    .o_dat    (ar_fifo_o_dat )
  );
  e603_subsys_gnrl_cdc_fifo # (
    .DP(ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (R_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_r(
    .o_clk   (icb_clk),
    .o_rst_n (icb_rst_n), 
    .i_clk   (async_axi_clk),
    .i_rst_n (async_axi_rst_n),
    .i_vld   (axi_rvalid),
    .i_rdy   (axi_rready),
    .i_dat   (r_fifo_i_dat ),
    .i_cdc_fifo_active(r_async_i_active),
    .o_cdc_fifo_active(r_async_o_active),
    .o_vld  (icb2axi_rvalid),
    .o_rdy  (icb2axi_rready),
    .o_dat  (r_fifo_o_dat )
  );
  wire axi2axi_async_i_active = ar_async_i_active | r_async_o_active ;
  wire axi2axi_async_o_active = ar_async_o_active | r_async_i_active ;
  assign icb2axi_read_async_icb_active = i_icb2axi_read_pend_active | axi2axi_async_i_active;
  assign icb2axi_read_async_axi_active = axi2axi_async_o_active;
  assign icb2axi_read_pend_active = icb2axi_read_async_icb_active;
endmodule
module e603_subsys_gnrl_ficb2axi_write_async_id # (
  parameter ID_W = 4,
  parameter SUPPORT_AWID_OOO = 0,
  parameter OUTS_CNT_W =2,
  parameter OUTS_FIFO_DP =4,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 1,
  parameter ASYNC_FIFO_DP = 6,
  parameter ASYNC_FIFO_DP_PTR_W = 3,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  output                        icb2axi_write_async_icb_active,
  output                        icb2axi_write_async_axi_active,
  output                        icb2axi_write_pend_active,
  input                         axi_awready,
  output                        axi_awvalid,
  output [AW-1:0]               axi_awaddr,
  output [7:0]                  axi_awlen,
  output [CMD_SIZE_W-1:0]                  axi_awsize,
  output [1:0]                  axi_awburst,
  output                        axi_awlock,
  output [3:0]                  axi_awcache,
  output [2:0]                  axi_awprot,
  output [CMD_UW-1:0]            axi_awuser, 
  output [ID_W-1:0]            axi_awid, 
  input                         axi_wready,
  output                        axi_wvalid,
  output [DW-1:0]               axi_wdata,
  output [DW/8-1:0]               axi_wstrb,
  output                        axi_wlast,
  output                         axi_bready,
  input                          axi_bvalid,
  input [RSP_UW-1:0]              axi_buser,
  input [ID_W-1:0]              axi_bid,
  input [1:0]                    axi_bresp,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [7:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input [ID_W-1:0]             icb_cmd_id,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]            icb_rsp_usr,
  output [ID_W-1:0]            icb_rsp_id,
  output                       icb_rsp_last,
  input  async_axi_clk,
  input  async_axi_rst_n,
  input  icb_clk,
  input  icb_rst_n
  );
  wire i_icb_reset_flag_r;
e603_subsys_gnrl_dffrs #(1) reset_flag_dffrs (1'b0, i_icb_reset_flag_r, icb_clk, icb_rst_n);// VPP_NO_REG_PARSE
  wire i_icb_cmd_valid;
  wire i_icb_cmd_ready;
  assign i_icb_cmd_valid = (~i_icb_reset_flag_r) & icb_cmd_valid;
  assign icb_cmd_ready   = (~i_icb_reset_flag_r) & i_icb_cmd_ready;
  wire aw_async_i_active;
  wire aw_async_o_active;
  wire w_async_i_active ;
  wire w_async_o_active ;
  wire b_async_o_active ;
  wire b_async_i_active ;
  wire axi2axi_async_i_active = aw_async_i_active | w_async_i_active | b_async_o_active ;
  wire axi2axi_async_o_active = aw_async_o_active | w_async_o_active | b_async_i_active ;
  wire                        icb2axi_awready;
  wire                        icb2axi_awvalid;
  wire [AW-1:0]               icb2axi_awaddr;
  wire [7:0]                  icb2axi_awlen;
  wire [CMD_SIZE_W-1:0]                  icb2axi_awsize;
  wire [1:0]                  icb2axi_awburst;
  wire                        icb2axi_awlock;
  wire [3:0]                  icb2axi_awcache;
  wire [2:0]                  icb2axi_awprot;
  wire [CMD_UW-1:0]           icb2axi_awuser;
  wire [ID_W-1:0]           icb2axi_awid;
  localparam AW_PACK_W = (AW+8+CMD_SIZE_W+2+1+4+3+CMD_UW+ID_W) 
                       ;
  wire [AW_PACK_W-1:0] aw_fifo_i_dat = {
                              icb2axi_awaddr,
                              icb2axi_awlen,
                              icb2axi_awsize,
                              icb2axi_awburst,
                              icb2axi_awlock,
                              icb2axi_awcache,
                              icb2axi_awprot,
                              icb2axi_awid, 
                              icb2axi_awuser 
                                 };
  wire [AW_PACK_W-1:0] aw_fifo_o_dat;
  assign {
                              axi_awaddr,
                              axi_awlen,
                              axi_awsize,
                              axi_awburst,
                              axi_awlock,
                              axi_awcache,
                              axi_awprot,
                              axi_awid,
                              axi_awuser
                                } = aw_fifo_o_dat;
  e603_subsys_gnrl_cdc_fifo # (
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (AW_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_aw(
    .i_clk   (icb_clk),
    .i_rst_n (icb_rst_n),
    .o_clk   (async_axi_clk),
    .o_rst_n (async_axi_rst_n),
    .i_vld    (icb2axi_awvalid),
    .i_rdy    (icb2axi_awready),
    .i_dat    (aw_fifo_i_dat),
    .i_cdc_fifo_active(aw_async_i_active),
    .o_cdc_fifo_active(aw_async_o_active),
    .o_vld    (axi_awvalid),
    .o_rdy    (axi_awready),
    .o_dat    (aw_fifo_o_dat )
  );
  wire                        icb2axi_wready;
  wire                        icb2axi_wvalid;
  wire [DW-1:0]               icb2axi_wdata;
  wire [DW/8-1:0]             icb2axi_wstrb;
  wire                        icb2axi_wlast;
  localparam W_PACK_W = (DW+(DW/8)+1);
  wire [W_PACK_W-1:0] w_fifo_i_dat = {
                              icb2axi_wdata,
                              icb2axi_wstrb,
                              icb2axi_wlast 
                                 };
  wire [W_PACK_W-1:0] w_fifo_o_dat;
  assign {
                              axi_wdata,
                              axi_wstrb,
                              axi_wlast 
                                } = w_fifo_o_dat;
  e603_subsys_gnrl_cdc_fifo # (
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (W_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_w(
    .i_clk   (icb_clk),
    .i_rst_n (icb_rst_n), 
    .o_clk   (async_axi_clk),
    .o_rst_n (async_axi_rst_n),
    .i_vld    (icb2axi_wvalid),
    .i_rdy    (icb2axi_wready),
    .i_dat    (w_fifo_i_dat),
    .i_cdc_fifo_active(w_async_i_active),
    .o_cdc_fifo_active(w_async_o_active),
    .o_vld    (axi_wvalid),
    .o_rdy    (axi_wready),
    .o_dat    (w_fifo_o_dat )
  );
  wire icb2axi_bvalid;
  wire icb2axi_bready;
  wire [RSP_UW-1:0] icb2axi_buser;
  wire [ID_W-1:0] icb2axi_bid;
  wire [1:0]        icb2axi_bresp;
  localparam B_PACK_W = (2+RSP_UW+ID_W);
  wire [B_PACK_W-1:0] b_fifo_i_dat = {
                                 axi_buser,
                                 axi_bid,
                                 axi_bresp 
                                 };
  wire [B_PACK_W-1:0] b_fifo_o_dat;
  assign {
                              icb2axi_buser,
                              icb2axi_bid,
                              icb2axi_bresp 
                                 } = b_fifo_o_dat;
  e603_subsys_gnrl_cdc_fifo # (
    .DP(ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (B_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_b(
    .o_clk   (icb_clk),
    .o_rst_n (icb_rst_n), 
    .i_clk   (async_axi_clk),
    .i_rst_n (async_axi_rst_n),
    .i_vld   (axi_bvalid),
    .i_rdy   (axi_bready),
    .i_dat   (b_fifo_i_dat ),
    .i_cdc_fifo_active(b_async_i_active),
    .o_cdc_fifo_active(b_async_o_active),
    .o_vld  (icb2axi_bvalid),
    .o_rdy  (icb2axi_bready),
    .o_dat  (b_fifo_o_dat )
  );
  wire i_icb2axi_write_pend_active;
 e603_subsys_gnrl_ficb2axi_write_id # (
            .ID_W (ID_W),
            .SUPPORT_AWID_OOO(SUPPORT_AWID_OOO),
            .AW (AW),
            .DW (DW),
            .RATIO_FIFO_DP(0),
            .OUTS_CNT_W  (OUTS_CNT_W ),
            .OUTS_FIFO_DP  (OUTS_FIFO_DP ),
            .CMD_UW (CMD_UW),
            .RSP_UW (RSP_UW)
   ) u_icb2axi_write(
            .icb2axi_write_pend_active(i_icb2axi_write_pend_active),
            .icb_cmd_valid   (i_icb_cmd_valid),
            .icb_cmd_ready   (i_icb_cmd_ready),
            .icb_cmd_addr    (icb_cmd_addr), 
            .icb_cmd_sel     (icb_cmd_sel), 
            .icb_cmd_xlen    (icb_cmd_xlen),
            .icb_cmd_xburst  (icb_cmd_xburst),
            .icb_cmd_modes   (icb_cmd_modes ),
            .icb_cmd_dmode   (icb_cmd_dmode ),
            .icb_cmd_attri   (icb_cmd_attri ),
            .icb_cmd_read    (icb_cmd_read), 
            .icb_cmd_wdata   (icb_cmd_wdata),
            .icb_cmd_wmask   (icb_cmd_wmask),
            .icb_cmd_beat    (icb_cmd_beat),
            .icb_cmd_lock    (icb_cmd_lock),
            .icb_cmd_excl    (icb_cmd_excl),
            .icb_cmd_size    (icb_cmd_size),
            .icb_cmd_usr     (icb_cmd_usr),
            .icb_cmd_id     (icb_cmd_id),
            .icb_rsp_valid   (icb_rsp_valid),
            .icb_rsp_ready   (icb_rsp_ready),
            .icb_rsp_rdata   (icb_rsp_rdata),
            .icb_rsp_usr     (icb_rsp_usr),
            .icb_rsp_err     (icb_rsp_err),
            .icb_rsp_excl_ok (icb_rsp_excl_ok),
            .icb_rsp_id (icb_rsp_id),
            .icb_rsp_last (icb_rsp_last),
            .axi_awready (icb2axi_awready ),
            .axi_awvalid (icb2axi_awvalid ),
            .axi_awaddr  (icb2axi_awaddr  ),
            .axi_awlen   (icb2axi_awlen   ),
            .axi_awsize  (icb2axi_awsize  ),
            .axi_awburst (icb2axi_awburst ),
            .axi_awlock  (icb2axi_awlock  ),
            .axi_awcache (icb2axi_awcache ),
            .axi_awprot  (icb2axi_awprot  ),
            .axi_awuser  (icb2axi_awuser  ),
            .axi_awid  (icb2axi_awid  ),
            .axi_wready  (icb2axi_wready  ),
            .axi_wvalid  (icb2axi_wvalid  ),
            .axi_wdata   (icb2axi_wdata   ),
            .axi_wstrb   (icb2axi_wstrb   ),
            .axi_wlast   (icb2axi_wlast   ),
            .axi_bready  (icb2axi_bready  ),
            .axi_bvalid  (icb2axi_bvalid  ),
            .axi_buser   (icb2axi_buser   ),
            .axi_bid   (icb2axi_bid   ),
            .axi_bresp   (icb2axi_bresp   ),
            .axi_bus_clk_en (1'b1),
            .icb_clk_en (1'b1),
            .clk   (icb_clk),
            .rst_n (icb_rst_n)
  );
  assign icb2axi_write_async_icb_active = i_icb2axi_write_pend_active | axi2axi_async_i_active;
  assign icb2axi_write_async_axi_active = axi2axi_async_o_active;
  assign icb2axi_write_pend_active = icb2axi_write_async_icb_active;
endmodule
`include "global.v"
module  e603_subsys_gnrl_axi2ficb_write_id # (
  parameter PAYLOAD_NORST = 0,
  parameter ALLOW_FIX_BURST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           axi_awready,
  input                            axi_awvalid,
  input [ID_W-1:0]        axi_awid,
  input [AW-1:0]      axi_awaddr,
  input [7:0]                      axi_awlen,
  input [CMD_SIZE_W-1:0]                      axi_awsize,
  input [1:0]                      axi_awburst,
  input                            axi_awlock,
  input [3:0]                      axi_awcache,
  input [2:0]                      axi_awprot,
  input [USR_W-1:0]          axi_awuser, 
  output                           axi_wready,
  input                            axi_wvalid,
  input [DW-1:0]           axi_wdata,
  input [MW-1:0]        axi_wstrb,
  input                            axi_wlast,
  input                            axi_bready,
  output                           axi_bvalid,
  output [USR_W-1:0]          axi_buser, 
  output [ID_W-1:0]       axi_bid,
  output [1:0]                     axi_bresp,
  output                           icb_wcmd_sel,
  output                           icb_wcmd_valid,
  input                            icb_wcmd_ready,
  output [AW-1:0]                  icb_wcmd_addr,
  output                           icb_wcmd_read, 
  output [DW-1:0]                  icb_wcmd_wdata,
  output [MW-1:0]                  icb_wcmd_wmask,
  output [1:0]                     icb_wcmd_beat,
  output                           icb_wcmd_lock,
  output                           icb_wcmd_excl,
  output [CMD_SIZE_W-1:0]         icb_wcmd_size,
  output [7:0]                     icb_wcmd_xlen,
  output [1:0]                     icb_wcmd_xburst,
  output [1:0]                     icb_wcmd_modes,
  output                           icb_wcmd_dmode,
  output [2:0]                     icb_wcmd_attri,
  output [USR_W-1:0]               icb_wcmd_usr,
  output [ID_W -1:0]               icb_wcmd_id,
  input                            icb_wrsp_valid,
  output                           icb_wrsp_ready,
  input                            icb_wrsp_err,
  input                            icb_wrsp_excl_ok,
  input  [USR_W-1:0]               icb_wrsp_usr,
  input [ID_W -1:0]                icb_wrsp_id,
  input                            axi_bus_clk_en,
  input                            icb_clk_en,
  output                           axi2icb_write_active,
  input  clk,
  input  rst_n
  );
  wire axi_awready_raw;
  wire axi_awvalid_raw;
  wire axi_wready_raw;
  wire axi_wvalid_raw;
  assign axi_awvalid_raw = (~reset_flag_r) & axi_awvalid    ;
  assign axi_awready     = (~reset_flag_r) & axi_awready_raw;
  assign axi_wvalid_raw  = (~reset_flag_r) & axi_wvalid    ;
  assign axi_wready      = (~reset_flag_r) & axi_wready_raw;
  assign icb_wcmd_lock = 1'b0;
    localparam AXI_AW_BUF_PACK = ID_W+AW+8+CMD_SIZE_W+2+1+3+4+USR_W;
    wire [AXI_AW_BUF_PACK-1:0] i_axi_aw_pack = {
                                             axi_awid    ,  
                                             axi_awaddr  ,
                                             axi_awlen   ,
                                             axi_awsize  ,
                                             axi_awburst ,
                                             axi_awlock  ,
                                             axi_awcache ,
                                             axi_awprot  ,
                                             axi_awuser   
                                            };
    wire [ID_W-1:0]    axi_buf_o_awid    ; 
    wire [AW-1:0]  axi_buf_o_awaddr  ; 
    wire [7:0]                  axi_buf_o_awlen   ; 
    wire [CMD_SIZE_W-1:0]                  axi_buf_o_awsize  ; 
    wire [1:0]                  axi_buf_o_awburst ; 
    wire                        axi_buf_o_awlock  ; 
    wire [3:0]                  axi_buf_o_awcache ; 
    wire [2:0]                  axi_buf_o_awprot  ; 
    wire [USR_W-1:0]      axi_buf_o_awuser  ; 
    wire [AXI_AW_BUF_PACK-1:0] o_axi_aw_pack ;
    assign  { 
              axi_buf_o_awid    , 
              axi_buf_o_awaddr  , 
              axi_buf_o_awlen   , 
              axi_buf_o_awsize  , 
              axi_buf_o_awburst , 
              axi_buf_o_awlock  , 
              axi_buf_o_awcache , 
              axi_buf_o_awprot  , 
              axi_buf_o_awuser    
            } = o_axi_aw_pack ;
    wire axi_buf_o_awvalid ;    
    wire axi_buf_o_awready ; 
    wire axi_o_awbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_AW_BUF_PACK)
    ) u_axi_aw_fifo(
    .i_clk_en(axi_bus_clk_en), 
    .i_vld(axi_awvalid_raw  ), 
    .i_rdy(axi_awready_raw  ), 
    .i_dat(i_axi_aw_pack),
    .o_clk_en(icb_clk_en),
    .o_vld(axi_buf_o_awvalid), 
    .o_rdy(axi_buf_o_awready), 
    .o_dat(o_axi_aw_pack    ),
    .o_fifo_active(axi_o_awbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
    localparam AXI_W_BUF_PACK = DW+MW+1;
    wire [AXI_W_BUF_PACK-1:0] i_axi_w_pack = {
                                             axi_wdata      , 
                                             axi_wstrb      , 
                                             axi_wlast        
                                            };
    wire [DW-1:0]       axi_buf_o_wdata  ; 
    wire [MW-1:0]    axi_buf_o_wstrb  ; 
    wire                        axi_buf_o_wlast  ; 
    wire [AXI_W_BUF_PACK-1:0] o_axi_w_pack ;
    assign  { 
              axi_buf_o_wdata  , 
              axi_buf_o_wstrb  , 
              axi_buf_o_wlast    
            } = o_axi_w_pack ;
    wire axi_buf_o_wvalid ;    
    wire axi_buf_o_wready ; 
    wire axi_o_wbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_W_BUF_PACK)
    ) u_axi_w_fifo(
    .i_clk_en(axi_bus_clk_en),
    .i_vld(axi_wvalid_raw  ), 
    .i_rdy(axi_wready_raw  ), 
    .i_dat(i_axi_w_pack),
    .o_clk_en(icb_clk_en),
    .o_vld(axi_buf_o_wvalid), 
    .o_rdy(axi_buf_o_wready), 
    .o_dat(o_axi_w_pack    ),
    .o_fifo_active(axi_o_wbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire axi_buf_o_awready_pos;
  wire axi_buf_o_awvalid_pos;
  wire write_id_fifo_rdy;
  assign axi_buf_o_awready     = write_id_fifo_rdy & axi_buf_o_awready_pos;
  assign axi_buf_o_awvalid_pos = write_id_fifo_rdy & axi_buf_o_awvalid    ;
  e603_subsys_gnrl_axi2ficb_aw_id # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W),
    .USR_W (USR_W)
  ) u_aw_axi2icb(
    .axi_awready  (axi_buf_o_awready_pos ),
    .axi_awvalid  (axi_buf_o_awvalid_pos & icb_clk_en ),
    .axi_awid     (axi_buf_o_awid    ),
    .axi_awaddr   (axi_buf_o_awaddr  ),
    .axi_awlen    (axi_buf_o_awlen   ),
    .axi_awsize   (axi_buf_o_awsize  ),
    .axi_awburst  (axi_buf_o_awburst ),
    .axi_awlock   (axi_buf_o_awlock  ),
    .axi_awcache  (axi_buf_o_awcache ),
    .axi_awprot   (axi_buf_o_awprot  ),
    .axi_awuser   (axi_buf_o_awuser),
    .axi_wready   (axi_buf_o_wready),
    .axi_wvalid   (axi_buf_o_wvalid & icb_clk_en),
    .axi_wdata    (axi_buf_o_wdata ),
    .axi_wstrb    (axi_buf_o_wstrb ),
    .axi_wlast    (axi_buf_o_wlast ),
    .icb_wcmd_sel (icb_wcmd_sel),
    .icb_wcmd_valid (icb_wcmd_valid),
    .icb_wcmd_ready (icb_wcmd_ready & icb_clk_en),
    .icb_wcmd_addr  (icb_wcmd_addr ), 
    .icb_wcmd_read  (icb_wcmd_read ), 
    .icb_wcmd_wdata (icb_wcmd_wdata),
    .icb_wcmd_wmask (icb_wcmd_wmask),
    .icb_wcmd_beat  (icb_wcmd_beat ),
    .icb_wcmd_lock  (              ), 
    .icb_wcmd_excl  (icb_wcmd_excl ),
    .icb_wcmd_size  (icb_wcmd_size ),
    .icb_wcmd_xlen    (icb_wcmd_xlen   ),
    .icb_wcmd_xburst  (icb_wcmd_xburst ),
    .icb_wcmd_modes   (icb_wcmd_modes  ),
    .icb_wcmd_dmode   (icb_wcmd_dmode  ),
    .icb_wcmd_attri   (icb_wcmd_attri  ),
    .icb_wcmd_usr   (icb_wcmd_usr  ), 
    .icb_wcmd_id    (icb_wcmd_id   ), 
    .clk (clk),
    .rst_n (rst_n)
  );
    localparam AXI_B_BUF_PACK = ID_W+2+USR_W;
    wire [USR_W-1:0]   axi_buf_i_buser    ; 
    wire [ID_W-1:0]    axi_buf_i_bid    ; 
    wire [1:0]                  axi_buf_i_bresp  ; 
    wire [AXI_B_BUF_PACK-1:0] i_axi_b_pack = {
                                             axi_buf_i_buser  ,  
                                             axi_buf_i_bid  ,  
                                             axi_buf_i_bresp        
                                            };
    wire [AXI_B_BUF_PACK-1:0] o_axi_b_pack ;
    assign  { 
              axi_buser    , 
              axi_bid    , 
              axi_bresp    
            } = o_axi_b_pack ;
    wire axi_buf_i_bvalid ;    
    wire axi_buf_i_bready ; 
    wire axi_o_bbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_B_BUF_PACK)
    ) u_axi_b_fifo(
    .i_clk_en(icb_clk_en),
    .i_vld(axi_buf_i_bvalid), 
    .i_rdy(axi_buf_i_bready), 
    .i_dat(i_axi_b_pack    ),
    .o_clk_en(axi_bus_clk_en),
    .o_vld(axi_bvalid  ), 
    .o_rdy(axi_bready  ), 
    .o_dat(o_axi_b_pack),
    .o_fifo_active(axi_o_bbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire write_id_fifo_active;
  wire [7:0] wrsp_xlen;
  wire  wrsp_burst;
  e603_subsys_gnrl_axi2ficb_b_id # (
    .USR_W (USR_W),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W)
  ) u_b_axi2icb(
    .icb_wrsp_ready   (icb_wrsp_ready  ),
    .icb_wrsp_valid   (icb_wrsp_valid  & icb_clk_en),
    .icb_wrsp_err     (icb_wrsp_err    ),
    .icb_wrsp_usr     (icb_wrsp_usr    ),
    .icb_wrsp_excl_ok (icb_wrsp_excl_ok),
    .icb_wrsp_id      (icb_wrsp_id   ), 
    .axi_bready       (axi_buf_i_bready & icb_clk_en),
    .axi_bvalid       (axi_buf_i_bvalid),
    .axi_bresp        (axi_buf_i_bresp ),
    .axi_buser        (axi_buf_i_buser ),
    .axi_bid          (axi_buf_i_bid   ), 
    .wrsp_xlen_vld  (write_id_fifo_active),
    .wrsp_xlen  (wrsp_xlen),
    .wrsp_burst (wrsp_burst),
    .clk (clk),
    .rst_n (rst_n)
  );
  wire wcmd_burst = (~(axi_buf_o_awlen == 8'b0)) ;
  wire [7:0] wcmd_xlen  = axi_buf_o_awlen;
  localparam WRSP_FIFO_PACK = 1+8+ID_W;
  e603_subsys_gnrl_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .CUT_READY (1),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
        .DW  (WRSP_FIFO_PACK)
  ) u_wrsp_fifo (
        .i_vld(axi_buf_o_awvalid && axi_buf_o_awready & icb_clk_en),
        .i_rdy(write_id_fifo_rdy),
        .i_dat({wcmd_burst,wcmd_xlen, axi_buf_o_awid}),
        .o_vld(write_id_fifo_active),
        .o_rdy(axi_buf_i_bvalid && axi_buf_i_bready & icb_clk_en ),  
        .o_dat({wrsp_burst,wrsp_xlen, 
                      axi_buf_i_bid
                      }),  
        .clk  (clk),
        .rst_n(rst_n)
  );
   assign axi2icb_write_active = axi_o_awbusy | axi_o_wbusy | axi_o_bbusy 
                               | write_id_fifo_active
                               ;
endmodule
module  e603_subsys_gnrl_axi2ficb_read_id # (
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           axi_arready,
  input                            axi_arvalid,
  input [ID_W-1:0]        axi_arid,
  input [AW-1:0]      axi_araddr,
  input [7:0]                      axi_arlen,
  input [CMD_SIZE_W-1:0]                      axi_arsize,
  input [1:0]                      axi_arburst,
  input                            axi_arlock,
  input [3:0]                      axi_arcache,
  input [2:0]                      axi_arprot,
  input [USR_W-1:0]          axi_aruser,
  input                            axi_rready,
  output                           axi_rvalid,
  output [ID_W-1:0]       axi_rid,
  output [DW-1:0]          axi_rdata,
  output [1:0]                     axi_rresp,
  output                           axi_rlast,
  output [USR_W-1:0]          axi_ruser,
  output                           icb_rcmd_sel ,
  output                           icb_rcmd_valid ,
  input                            icb_rcmd_ready ,
  output [AW-1:0]                  icb_rcmd_addr  ,
  output                           icb_rcmd_read  ,
  output [DW-1:0]                  icb_rcmd_wdata ,
  output [MW-1:0]                  icb_rcmd_wmask ,
  output [1:0]                     icb_rcmd_beat  ,
  output                           icb_rcmd_excl  ,             
  output [CMD_SIZE_W-1:0]         icb_rcmd_size  ,
  output [7:0]                     icb_rcmd_xlen,
  output [1:0]                     icb_rcmd_xburst,
  output [1:0]                     icb_rcmd_modes,
  output                           icb_rcmd_dmode,
  output [2:0]                     icb_rcmd_attri,
  output [USR_W-1:0]               icb_rcmd_usr   ,
  output [ID_W -1:0]               icb_rcmd_id   ,
  output                           icb_rrsp_ready  , 
  input                            icb_rrsp_valid  , 
  input [DW-1:0]                   icb_rrsp_rdata  , 
  input                            icb_rrsp_err    , 
  input                            icb_rrsp_excl_ok, 
  input [USR_W-1:0]                icb_rrsp_usr   ,
  input [ID_W -1:0]                icb_rrsp_id   ,
  input                            icb_rrsp_last,
  input                            axi_bus_clk_en,
  input                            icb_clk_en,
  output                           axi2icb_read_active,
  input clk  ,
  input rst_n  
  );
  wire axi_arvalid_raw;
  wire axi_arready_raw;
  assign axi_arvalid_raw = (~reset_flag_r) & axi_arvalid;
  assign axi_arready     = (~reset_flag_r) & axi_arready_raw;
    localparam AXI_AR_BUF_PACK = ID_W+AW+8+CMD_SIZE_W+2+1+3+4+USR_W;
    wire [AXI_AR_BUF_PACK-1:0] i_axi_ar_pack = {
                                             axi_arid    ,  
                                             axi_araddr  ,
                                             axi_arlen   ,
                                             axi_arsize  ,
                                             axi_arburst ,
                                             axi_arlock  ,
                                             axi_arcache ,
                                             axi_arprot  ,
                                             axi_aruser   
                                            };
    wire [ID_W-1:0]    axi_buf_o_arid    ; 
    wire [AW-1:0]  axi_buf_o_araddr  ; 
    wire [7:0]                  axi_buf_o_arlen   ; 
    wire [CMD_SIZE_W-1:0]                  axi_buf_o_arsize  ; 
    wire [1:0]                  axi_buf_o_arburst ; 
    wire                        axi_buf_o_arlock  ; 
    wire [3:0]                  axi_buf_o_arcache ; 
    wire [2:0]                  axi_buf_o_arprot  ; 
    wire [USR_W-1:0]      axi_buf_o_aruser  ; 
    wire [AXI_AR_BUF_PACK-1:0] o_axi_ar_pack ;
    assign  { 
              axi_buf_o_arid    , 
              axi_buf_o_araddr  , 
              axi_buf_o_arlen   , 
              axi_buf_o_arsize  , 
              axi_buf_o_arburst , 
              axi_buf_o_arlock  , 
              axi_buf_o_arcache , 
              axi_buf_o_arprot  , 
              axi_buf_o_aruser    
            } = o_axi_ar_pack ;
    wire axi_buf_o_arvalid ;    
    wire axi_buf_o_arready ; 
    wire axi_o_arbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_AR_BUF_PACK)
    ) u_axi_ar_fifo(
    .i_clk_en(axi_bus_clk_en), 
    .i_vld(axi_arvalid_raw      ), 
    .i_rdy(axi_arready_raw      ), 
    .i_dat(i_axi_ar_pack    ),
    .o_clk_en(icb_clk_en), 
    .o_vld(axi_buf_o_arvalid), 
    .o_rdy(axi_buf_o_arready), 
    .o_dat(o_axi_ar_pack    ),
    .o_fifo_active(axi_o_arbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire axi_buf_o_arready_pos;
  wire axi_buf_o_arvalid_pos;
  wire read_id_fifo_rdy;
  assign axi_buf_o_arready     = read_id_fifo_rdy & axi_buf_o_arready_pos;
  assign axi_buf_o_arvalid_pos = read_id_fifo_rdy & axi_buf_o_arvalid;
  e603_subsys_gnrl_axi2ficb_ar_id # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W),
    .USR_W (USR_W)  
  ) u_ar_axi2icb(
     .axi_arready  (axi_buf_o_arready_pos ),
     .axi_arvalid  (axi_buf_o_arvalid_pos & icb_clk_en ),
     .axi_arid     (axi_buf_o_arid    ),
     .axi_araddr   (axi_buf_o_araddr  ),
     .axi_arlen    (axi_buf_o_arlen   ),
     .axi_arsize   (axi_buf_o_arsize  ),
     .axi_arburst  (axi_buf_o_arburst ),
     .axi_arlock   (axi_buf_o_arlock  ),
     .axi_arcache  (axi_buf_o_arcache ),
     .axi_arprot   (axi_buf_o_arprot  ),
     .axi_aruser   (axi_buf_o_aruser), 
     .icb_rcmd_sel   (icb_rcmd_sel),
     .icb_rcmd_valid (icb_rcmd_valid),
     .icb_rcmd_ready (icb_rcmd_ready & icb_clk_en),
     .icb_rcmd_addr  (icb_rcmd_addr ), 
     .icb_rcmd_read  (icb_rcmd_read ), 
     .icb_rcmd_wdata (icb_rcmd_wdata),
     .icb_rcmd_wmask (icb_rcmd_wmask),
     .icb_rcmd_beat  (icb_rcmd_beat ),
     .icb_rcmd_lock  (              ), 
     .icb_rcmd_excl  (icb_rcmd_excl ),
     .icb_rcmd_size  (icb_rcmd_size ),
     .icb_rcmd_xlen    (icb_rcmd_xlen   ),
     .icb_rcmd_xburst  (icb_rcmd_xburst ),
     .icb_rcmd_modes   (icb_rcmd_modes  ),
     .icb_rcmd_dmode   (icb_rcmd_dmode  ),
     .icb_rcmd_attri   (icb_rcmd_attri  ),
     .icb_rcmd_usr   (icb_rcmd_usr  ),
     .icb_rcmd_id    (icb_rcmd_id   ),
     .clk   (clk),
     .rst_n (rst_n)
  );
    localparam AXI_R_BUF_PACK = USR_W+ID_W+DW+2+1;
    wire [USR_W-1:0]    axi_buf_i_ruser    ; 
    wire [ID_W-1:0]    axi_buf_i_rid    ; 
    wire [DW-1:0]       axi_buf_i_rdata  ; 
    wire [1:0]                  axi_buf_i_rresp  ; 
    wire                        axi_buf_i_rlast  ; 
    wire [AXI_R_BUF_PACK-1:0] i_axi_r_pack = {
                                             axi_buf_i_ruser    ,
                                             axi_buf_i_rid    ,
                                             axi_buf_i_rdata  ,
                                             axi_buf_i_rresp  ,
                                             axi_buf_i_rlast   
                                            };
    wire [AXI_R_BUF_PACK-1:0] o_axi_r_pack ;
    assign  { 
              axi_ruser        ,  
              axi_rid        ,  
              axi_rdata      ,  
              axi_rresp      ,  
              axi_rlast         
            } = o_axi_r_pack ;
    wire axi_buf_i_rvalid ;    
    wire axi_buf_i_rready ; 
    wire axi_o_rbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_R_BUF_PACK)
    ) u_axi_r_fifo(
    .i_clk_en(icb_clk_en),
    .i_vld(axi_buf_i_rvalid), 
    .i_rdy(axi_buf_i_rready), 
    .i_dat(i_axi_r_pack    ),
    .o_clk_en(axi_bus_clk_en),
    .o_vld(axi_rvalid  ), 
    .o_rdy(axi_rready  ), 
    .o_dat(o_axi_r_pack),
    .o_fifo_active(axi_o_rbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire read_id_fifo_active;
  e603_subsys_gnrl_axi2ficb_r_id # (
    .USR_W (USR_W),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W)
  ) u_axi2icb_r(
    .icb_rrsp_ready   (icb_rrsp_ready  ),
    .icb_rrsp_valid   (icb_rrsp_valid  & icb_clk_en  ),
    .icb_rrsp_rdata   (icb_rrsp_rdata  ),
    .icb_rrsp_usr     (icb_rrsp_usr    ),
    .icb_rrsp_err     (icb_rrsp_err    ),
    .icb_rrsp_excl_ok (icb_rrsp_excl_ok),
     .icb_rrsp_id     (icb_rrsp_id   ),
     .icb_rrsp_last   (icb_rrsp_last ),
    .axi_rready       (axi_buf_i_rready & icb_clk_en),
    .axi_rvalid       (axi_buf_i_rvalid),
    .axi_rid          (axi_buf_i_rid   ),
    .axi_ruser        (axi_buf_i_ruser ),
    .axi_rdata        (axi_buf_i_rdata ),
    .axi_rresp        (axi_buf_i_rresp ),
    .axi_rlast        (axi_buf_i_rlast ),
    .clk   (clk          ),
    .rst_n (rst_n)
  );
  localparam RRSP_FIFO_PACK = 1+8+ID_W;
  e603_subsys_gnrl_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .CUT_READY (1),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM), 
        .DW  (1)
  ) u_rrsp_fifo (
        .i_vld(axi_buf_o_arvalid && axi_buf_o_arready  & icb_clk_en), 
        .i_rdy(read_id_fifo_rdy),
        .o_vld(read_id_fifo_active),
        .o_rdy(axi_buf_i_rvalid && axi_buf_i_rready && axi_buf_i_rlast  & icb_clk_en ),  
        .i_dat(1'b0),
        .o_dat(),  
        .clk  (clk),
        .rst_n(rst_n)
  );
  assign axi2icb_read_active = axi_o_arbusy | axi_o_rbusy 
                             | read_id_fifo_active
                             ;
endmodule
module  e603_subsys_gnrl_axi2ficb_ar_id # (
  parameter PAYLOAD_NORST = 0,
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ID_W = 4, 
  parameter USR_W = 1
) (
  output                         axi_arready,
  input                          axi_arvalid,
  input [ID_W-1:0]               axi_arid,
  input [AW-1:0]                 axi_araddr,
  input [7:0]                    axi_arlen,
  input [CMD_SIZE_W-1:0]                    axi_arsize,
  input [1:0]                    axi_arburst,
  input                          axi_arlock,
  input [3:0]                    axi_arcache,
  input [2:0]                    axi_arprot,
  input [USR_W-1:0]              axi_aruser,
  output                         icb_rcmd_valid,
  input                          icb_rcmd_ready,
  output [AW-1:0]                icb_rcmd_addr, 
  output                         icb_rcmd_read, 
  output [DW-1:0]                icb_rcmd_wdata,
  output [MW-1:0]                icb_rcmd_wmask,
  output [1:0]                   icb_rcmd_beat,
  output                         icb_rcmd_lock,
  output                         icb_rcmd_excl,
  output [CMD_SIZE_W-1:0]       icb_rcmd_size,
  output [USR_W-1:0]             icb_rcmd_usr,
  output                         icb_rcmd_sel,
  output [7:0]                   icb_rcmd_xlen,
  output [1:0]                   icb_rcmd_xburst,
  output [1:0]                   icb_rcmd_modes,
  output                         icb_rcmd_dmode,
  output [2:0]                   icb_rcmd_attri,
  output[ID_W-1:0]               icb_rcmd_id,
  input                         clk,
  input                         rst_n
  );
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_nxt;
  wire       burst_cnt_ena;
  wire       rcmd_burst;
  wire       rcmd_burst_r;
  wire axi_arlock_buf;
  wire [CMD_SIZE_W-1:0] axi_arsize_buf;
  wire [1:0] axi_arburst_buf;
  wire [7:0] axi_arlen_buf;
  wire [2:0] axi_arprot_buf ;
  wire [3:0] axi_arcache_buf;
  wire [USR_W-1:0] axi_aruser_buf;
  wire [ID_W-1:0] axi_arid_buf;
  wire [AW-1:0] axi_araddr_buf;
  wire buf_wr_en;
  assign rcmd_burst = axi_arvalid  & (~(axi_arlen == 8'b0)) ;
  wire burst_first = (burst_cnt_r == 8'b0);
  assign rcmd_burst_r = ~burst_first;
  assign burst_cnt_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_last = (burst_cnt_r == axi_arlen_buf) & (~burst_first);
  assign burst_cnt_ena = (rcmd_burst || rcmd_burst_r) && icb_rcmd_valid && icb_rcmd_ready;
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign buf_wr_en = rcmd_burst && icb_rcmd_valid && icb_rcmd_ready && burst_first;
  generate
  if(PAYLOAD_NORST == 1) begin: payload_norst 
e603_subsys_gnrl_dffl  #(1) arlock_dffl  ( buf_wr_en, axi_arlock, axi_arlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(CMD_SIZE_W) arsize_dffl  ( buf_wr_en, axi_arsize, axi_arsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(8) arlen_dffl  ( buf_wr_en, axi_arlen, axi_arlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2) arburst_dffl  ( buf_wr_en, axi_arburst, axi_arburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(USR_W) aruser_dffl  ( buf_wr_en, axi_aruser, axi_aruser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(3) arprot_dffl   ( buf_wr_en, axi_arprot,  axi_arprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(4) arcache_dffl  ( buf_wr_en, axi_arcache, axi_arcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(ID_W) arid_dffl  ( buf_wr_en, axi_arid, axi_arid_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: payload_rst
e603_subsys_gnrl_dfflr #(1) arlock_dfflr ( buf_wr_en, axi_arlock, axi_arlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(CMD_SIZE_W) arsize_dfflr ( buf_wr_en, axi_arsize, axi_arsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(8) arlen_dfflr ( buf_wr_en, axi_arlen, axi_arlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(2) arburst_dfflr ( buf_wr_en, axi_arburst, axi_arburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(USR_W) aruser_dfflr ( buf_wr_en, axi_aruser, axi_aruser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(3) arprot_dfflr  ( buf_wr_en, axi_arprot,  axi_arprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(4) arcache_dfflr ( buf_wr_en, axi_arcache, axi_arcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(ID_W) arid_dfflr ( buf_wr_en, axi_arid, axi_arid_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  assign axi_arready   = icb_rcmd_ready && (!rcmd_burst_r);
  assign icb_rcmd_valid   = axi_arvalid  || rcmd_burst_r;
  wire icb_rcmd_read_tmp    = 1'b1; 
  assign icb_rcmd_read = icb_rcmd_read_tmp;
  assign icb_rcmd_wdata   = {DW{1'b0}};
  assign icb_rcmd_wmask   = {MW{1'b0}};
  wire icb_rcmd_lock_tmp    = 1'b0; 
  assign icb_rcmd_lock    = icb_rcmd_lock_tmp;
  wire icb_rcmd_excl_tmp    = rcmd_burst_r ? axi_arlock_buf : axi_arlock;
  assign icb_rcmd_excl = icb_rcmd_excl_tmp;
  wire [CMD_SIZE_W-1:0] icb_rcmd_size_tmp;
  assign icb_rcmd_size_tmp    = rcmd_burst_r ? axi_arsize_buf[CMD_SIZE_W-1:0] : axi_arsize[CMD_SIZE_W-1:0];
  assign icb_rcmd_size = icb_rcmd_size_tmp;
  wire icb_rcmd_fxed;
  wire icb_rcmd_incr;
  wire icb_rcmd_wrap;
  wire axi_araddr_ena = burst_cnt_ena;
  wire [AW-1:0] icb_rcmd_addr_mask = ({AW{1'b1}} << icb_rcmd_size);
  wire [AW-1:0] icb_rcmd_addr_algned = (icb_rcmd_addr_mask & icb_rcmd_addr);
  wire [12-1:0] axi_araddr_incr_size = (icb_rcmd_addr_algned[11:0] + (12'b1 << icb_rcmd_size));
  wire [12-1:0] axi_araddr_wrap_mask = ((~{8'b0,icb_rcmd_xlen[3:0]}) << icb_rcmd_size);
  wire [12-1:0] axi_araddr_incr_wrap = (axi_araddr_incr_size & (~axi_araddr_wrap_mask)) | (icb_rcmd_addr[11:0] & axi_araddr_wrap_mask);
  wire [AW-1:0] axi_araddr_nxt = icb_rcmd_fxed ? icb_rcmd_addr : 
                                 icb_rcmd_wrap ? {icb_rcmd_addr[AW-1:12],axi_araddr_incr_wrap} :
                                                 {icb_rcmd_addr[AW-1:12],axi_araddr_incr_size};
  generate
  if(PAYLOAD_NORST == 1) begin: araddr_payload_norst 
e603_subsys_gnrl_dffl  #(AW) araddr_dffl  ( axi_araddr_ena, axi_araddr_nxt, axi_araddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: araddr_payload_rst
e603_subsys_gnrl_dfflr #(AW) araddr_dfflr ( axi_araddr_ena, axi_araddr_nxt, axi_araddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  wire icb_rcmd_xlen_eq3  = (icb_rcmd_xlen == 8'd3) ;
  wire icb_rcmd_xlen_eq7  = (icb_rcmd_xlen == 8'd7) ;
  wire icb_rcmd_xlen_eq15 = (icb_rcmd_xlen == 8'd15);
  assign icb_rcmd_fxed = (icb_rcmd_xburst == 2'b00);
  assign icb_rcmd_incr = (icb_rcmd_xburst == 2'b01);
  assign icb_rcmd_wrap = (icb_rcmd_xburst == 2'b10);
  wire icb_rcmd_xburst_fixed;
  wire [1:0] icb_rcmd_beat_tmp;
  assign icb_rcmd_beat_tmp  = icb_rcmd_xburst_fixed          ? 2'b00 :
                          ( rcmd_burst && !rcmd_burst_r) ? 2'b01 : 
                          (burst_last)                   ? 2'b10 :
                                                           2'b00 ;
  assign icb_rcmd_beat = icb_rcmd_beat_tmp;
  wire [AW-1:0] icb_rcmd_addr_raw; 
  assign icb_rcmd_addr_raw  = (!rcmd_burst_r) ? axi_araddr :
                          axi_araddr_buf ; 
  assign icb_rcmd_usr   = rcmd_burst_r ? axi_aruser_buf : axi_aruser;
  wire [ID_W-1:0] icb_rcmd_id_tmp;
  assign icb_rcmd_id_tmp    = rcmd_burst_r ? axi_arid_buf   : axi_arid;
  assign icb_rcmd_id = icb_rcmd_id_tmp; 
  wire [2:0] icb_rcmd_arprot  = rcmd_burst_r ? axi_arprot_buf  : axi_arprot;
  wire [3:0] icb_rcmd_arcache = rcmd_burst_r ? axi_arcache_buf : axi_arcache;
  wire [7:0] icb_rcmd_arlen   = rcmd_burst_r ? axi_arlen_buf   : axi_arlen;
  wire [AW-1:0] icb_rcmd_addr_tmp;
  assign icb_rcmd_addr_tmp  = icb_rcmd_addr_raw;
  assign icb_rcmd_addr = icb_rcmd_addr_tmp; 
  wire icb_rcmd_nonalloc = (icb_rcmd_arcache == 4'b1011);
  wire icb_rcmd_device = icb_rcmd_nonalloc | (icb_rcmd_arcache == 4'b0000) | (icb_rcmd_arcache == 4'b0001);
  wire icb_rcmd_cacheb = (icb_rcmd_arcache == 4'b1111) | (icb_rcmd_arcache == 4'b0111) | (icb_rcmd_arcache == 4'b1011);
  wire icb_rcmd_nc     = icb_rcmd_nonalloc | ((~icb_rcmd_device) & (~icb_rcmd_cacheb));
  wire icb_rcmd_mmode = icb_rcmd_arprot[0];
  wire icb_rcmd_hmode = 1'b0;
  wire icb_rcmd_smode = 1'b0;
  wire icb_rcmd_ifu   = icb_rcmd_arprot[2];
  assign icb_rcmd_sel  = icb_rcmd_valid;
  wire [1:0] icb_rcmd_modes_tmp;
  assign icb_rcmd_modes_tmp = icb_rcmd_mmode ? 2'd0 : icb_rcmd_hmode ? 2'd1 : icb_rcmd_smode ? 2'd2 : 2'd3;
  assign icb_rcmd_modes = icb_rcmd_modes_tmp;
  wire icb_rcmd_dmode_tmp = 1'b0;
  assign icb_rcmd_dmode = icb_rcmd_dmode_tmp;
  wire [2:0] icb_rcmd_attri_tmp;
  assign icb_rcmd_attri_tmp[0] = icb_rcmd_ifu   ;
  assign icb_rcmd_attri_tmp[1] = icb_rcmd_device;
  assign icb_rcmd_attri_tmp[2] = icb_rcmd_nc    ;
  assign icb_rcmd_attri = icb_rcmd_attri_tmp;
  wire [7:0] icb_rcmd_xlen_tmp;
  assign icb_rcmd_xlen_tmp = icb_rcmd_xburst_fixed ? 8'd0 : icb_rcmd_arlen;
  assign icb_rcmd_xlen = icb_rcmd_xlen_tmp;
  generate 
      if(ALLOW_FIX_BURST == 1) begin: allow_fix_burst_gen
  assign icb_rcmd_xburst_fixed = 1'b0;
      end
      else begin: disallow_fix_burst_gen
  assign icb_rcmd_xburst_fixed = (icb_rcmd_xburst == 2'b00);
      end
  endgenerate
  wire [1:0] icb_rcmd_xburst_tmp; 
  assign icb_rcmd_xburst_tmp = rcmd_burst_r ? axi_arburst_buf : axi_arburst;
  assign icb_rcmd_xburst = icb_rcmd_xburst_tmp;
endmodule
module  e603_subsys_gnrl_axi2ficb_aw_id # (
  parameter PAYLOAD_NORST = 0,
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  output                         axi_awready,
  input                          axi_awvalid,
  input [ID_W-1:0]               axi_awid,
  input [AW-1:0]                 axi_awaddr,
  input [7:0]                    axi_awlen,
  input [CMD_SIZE_W-1:0]                    axi_awsize,
  input [1:0]                    axi_awburst,
  input                          axi_awlock,
  input [3:0]                    axi_awcache,
  input [2:0]                    axi_awprot,
  input [USR_W-1:0]              axi_awuser,
  output                         axi_wready,
  input                          axi_wvalid,
  input [DW-1:0]                 axi_wdata,
  input [MW-1:0]                 axi_wstrb,
  input                          axi_wlast,
  output                         icb_wcmd_valid,
  input                          icb_wcmd_ready,
  output [AW-1:0]                icb_wcmd_addr, 
  output                         icb_wcmd_read, 
  output [DW-1:0]                icb_wcmd_wdata,
  output [MW-1:0]                icb_wcmd_wmask,
  output [1:0]                   icb_wcmd_beat,
  output                         icb_wcmd_lock,
  output                         icb_wcmd_excl,
  output [CMD_SIZE_W-1:0]       icb_wcmd_size,
  output [USR_W-1:0]             icb_wcmd_usr,
  output                         icb_wcmd_sel,
  output [7:0]                   icb_wcmd_xlen,
  output [1:0]                   icb_wcmd_xburst,
  output [1:0]                   icb_wcmd_modes,
  output                         icb_wcmd_dmode,
  output [2:0]                   icb_wcmd_attri,
  output [ID_W-1:0]              icb_wcmd_id,
  input                         clk,
  input                         rst_n
  );
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_nxt;
  wire       burst_cnt_ena;
  wire       wcmd_burst;
  wire       wcmd_burst_r;
  wire axi_awlock_buf;
  wire [CMD_SIZE_W-1:0] axi_awsize_buf;
  wire [1:0] axi_awburst_buf;
  wire [7:0] axi_awlen_buf;
  wire [USR_W-1:0] axi_awuser_buf;
  wire [ID_W-1:0] axi_awid_buf;
  wire [AW-1:0] axi_awaddr_buf;
  wire [2:0] axi_awprot_buf ;
  wire [3:0] axi_awcache_buf;
  wire buf_wr_en;
  assign wcmd_burst = axi_awvalid  & (~(axi_awlen == 8'b0)) ;
  wire burst_first = (burst_cnt_r == 8'b0);
  assign wcmd_burst_r = ~burst_first;
  assign burst_cnt_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_last = (burst_cnt_r == axi_awlen_buf)& (~burst_first);
  assign burst_cnt_ena = (wcmd_burst || wcmd_burst_r) && icb_wcmd_valid && icb_wcmd_ready;
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign buf_wr_en = wcmd_burst && icb_wcmd_valid && icb_wcmd_ready && burst_first;
  generate
  if(PAYLOAD_NORST == 1) begin: payload_norst 
e603_subsys_gnrl_dffl  #(1) awlock_dffl  ( buf_wr_en, axi_awlock, axi_awlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(CMD_SIZE_W) awsize_dffl  ( buf_wr_en, axi_awsize, axi_awsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(8) awlen_dffl  ( buf_wr_en, axi_awlen, axi_awlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2) awburst_dffl  ( buf_wr_en, axi_awburst, axi_awburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(USR_W) awuser_dffl  ( buf_wr_en, axi_awuser, axi_awuser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(ID_W) awid_dffl  ( buf_wr_en, axi_awid, axi_awid_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(3) awprot_dffl   ( buf_wr_en, axi_awprot,  axi_awprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(4) awcache_dffl  ( buf_wr_en, axi_awcache, axi_awcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: payload_rst
e603_subsys_gnrl_dfflr #(1) awlock_dfflr ( buf_wr_en, axi_awlock, axi_awlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(CMD_SIZE_W) awsize_dfflr ( buf_wr_en, axi_awsize, axi_awsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(8) awlen_dfflr ( buf_wr_en, axi_awlen, axi_awlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(2) awburst_dfflr ( buf_wr_en, axi_awburst, axi_awburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(USR_W) awuser_dfflr ( buf_wr_en, axi_awuser, axi_awuser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(ID_W) awid_dfflr ( buf_wr_en, axi_awid, axi_awid_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(3) awprot_dfflr  ( buf_wr_en, axi_awprot,  axi_awprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(4) awcache_dfflr ( buf_wr_en, axi_awcache, axi_awcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  wire icb_wcmd_read_tmp; 
  assign icb_wcmd_read_tmp    = 1'b0; 
  assign icb_wcmd_read = icb_wcmd_read_tmp;
  wire [DW-1:0] icb_wcmd_wdata_tmp;
  wire [MW-1:0] icb_wcmd_wmask_tmp;
  assign icb_wcmd_wdata_tmp   = axi_wdata;
  assign icb_wcmd_wmask_tmp   = axi_wstrb;
  assign icb_wcmd_wdata = icb_wcmd_wdata_tmp;
  assign icb_wcmd_wmask = icb_wcmd_wmask_tmp;
  wire [CMD_SIZE_W-1:0] icb_wcmd_size_tmp;
  wire icb_wcmd_lock_tmp    = 1'b0;
  assign icb_wcmd_lock = icb_wcmd_lock_tmp;
  wire icb_wcmd_excl_tmp    = wcmd_burst_r ? axi_awlock_buf : axi_awlock;
  assign icb_wcmd_excl = icb_wcmd_excl_tmp;
  assign icb_wcmd_size_tmp    = wcmd_burst_r ? axi_awsize_buf[CMD_SIZE_W-1:0] : axi_awsize[CMD_SIZE_W-1:0];
  assign icb_wcmd_size    = icb_wcmd_size_tmp;
  assign axi_awready   = icb_wcmd_ready && (!wcmd_burst_r) && axi_wvalid;
  assign axi_wready    = icb_wcmd_ready && (wcmd_burst_r || axi_awvalid);
  assign icb_wcmd_valid   = (axi_awvalid || wcmd_burst_r) && axi_wvalid ;
  wire icb_wcmd_fxed;
  wire icb_wcmd_incr;
  wire icb_wcmd_wrap;
  wire axi_awaddr_ena = burst_cnt_ena;
  wire [AW-1:0] icb_wcmd_addr_mask = ({AW{1'b1}} << icb_wcmd_size);
  wire [AW-1:0] icb_wcmd_addr_algned = (icb_wcmd_addr_mask & icb_wcmd_addr);
  wire [12-1:0] axi_awaddr_incr_size = (icb_wcmd_addr_algned[11:0] + (12'b1 << icb_wcmd_size));
  wire [12-1:0] axi_awaddr_wrap_mask = ((~{8'b0,icb_wcmd_xlen[3:0]}) << icb_wcmd_size);
  wire [12-1:0] axi_awaddr_incr_wrap = (axi_awaddr_incr_size & (~axi_awaddr_wrap_mask)) | (icb_wcmd_addr[11:0] & axi_awaddr_wrap_mask);
  wire [AW-1:0] axi_awaddr_nxt = icb_wcmd_fxed ? icb_wcmd_addr : 
                                 icb_wcmd_wrap ? {icb_wcmd_addr[AW-1:12],axi_awaddr_incr_wrap} :
                                                 {icb_wcmd_addr[AW-1:12],axi_awaddr_incr_size};
    generate
  if(PAYLOAD_NORST == 1) begin: awaddr_payload_norst 
e603_subsys_gnrl_dffl  #(AW) awaddr_dffl  ( axi_awaddr_ena, axi_awaddr_nxt, axi_awaddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: awaddr_payload_rst
e603_subsys_gnrl_dfflr #(AW) awaddr_dfflr ( axi_awaddr_ena, axi_awaddr_nxt, axi_awaddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  wire icb_wcmd_xlen_eq3  = (icb_wcmd_xlen == 8'd3) ;
  wire icb_wcmd_xlen_eq7  = (icb_wcmd_xlen == 8'd7) ;
  wire icb_wcmd_xlen_eq15 = (icb_wcmd_xlen == 8'd15);
  assign icb_wcmd_fxed = (icb_wcmd_xburst == 2'b00);
  assign icb_wcmd_incr = (icb_wcmd_xburst == 2'b01);
  assign icb_wcmd_wrap = (icb_wcmd_xburst == 2'b10);
  wire icb_wcmd_xburst_fixed;
  wire [1:0] icb_wcmd_beat_tmp;
  assign icb_wcmd_beat_tmp  = icb_wcmd_xburst_fixed          ? 
                                        2'b00 :
                          ( wcmd_burst && !wcmd_burst_r) ? 2'b01 : 
                          (burst_last)                   ? 2'b10 :
                                                           2'b00 ;
  assign icb_wcmd_beat  = icb_wcmd_beat_tmp;
  wire [AW-1:0] icb_wcmd_addr_raw; 
  assign icb_wcmd_addr_raw  = (!wcmd_burst_r) ? axi_awaddr :
                          axi_awaddr_buf ; 
  assign icb_wcmd_usr   = wcmd_burst_r ? axi_awuser_buf : axi_awuser;
  wire [ID_W-1:0] icb_wcmd_id_tmp;
  assign icb_wcmd_id_tmp    = {ID_W{1'b0}};
  assign icb_wcmd_id = icb_wcmd_id_tmp; 
  wire [2:0] icb_wcmd_awprot  = wcmd_burst_r ? axi_awprot_buf  : axi_awprot;
  wire [3:0] icb_wcmd_awcache = wcmd_burst_r ? axi_awcache_buf : axi_awcache;
  wire [7:0] icb_wcmd_awlen   = wcmd_burst_r ? axi_awlen_buf   : axi_awlen;
  wire [AW-1:0] icb_wcmd_addr_tmp;
  assign icb_wcmd_addr_tmp  = icb_wcmd_addr_raw;
  assign icb_wcmd_addr = icb_wcmd_addr_tmp;  
  wire icb_wcmd_nonalloc = (icb_wcmd_awcache == 4'b0111);
  wire icb_wcmd_device = icb_wcmd_nonalloc | (icb_wcmd_awcache == 4'b0000) | (icb_wcmd_awcache == 4'b0001);
  wire icb_wcmd_cacheb = (icb_wcmd_awcache == 4'b1111) | (icb_wcmd_awcache == 4'b0111) | (icb_wcmd_awcache == 4'b1011);
  wire icb_wcmd_nc     = icb_wcmd_nonalloc | ((~icb_wcmd_device) & (~icb_wcmd_cacheb));
  wire icb_wcmd_mmode = icb_wcmd_awprot[0];
  wire icb_wcmd_hmode = 1'b0;
  wire icb_wcmd_smode = 1'b0;
  wire icb_wcmd_ifu   = icb_wcmd_awprot[2];
  assign icb_wcmd_sel  = icb_wcmd_valid;
  wire [1:0] icb_wcmd_modes_tmp = icb_wcmd_mmode ? 2'd0 : icb_wcmd_hmode ? 2'd1 : icb_wcmd_smode ? 2'd2 : 2'd3;
  assign icb_wcmd_modes = icb_wcmd_modes_tmp;
  wire icb_wcmd_dmode_tmp = 1'b0;
  wire [2:0] icb_wcmd_attri_tmp;
  assign icb_wcmd_dmode = icb_wcmd_dmode_tmp;
  assign icb_wcmd_attri_tmp[0] = icb_wcmd_ifu   ;
  assign icb_wcmd_attri_tmp[1] = icb_wcmd_device;
  assign icb_wcmd_attri_tmp[2] = icb_wcmd_nc    ;
  assign icb_wcmd_attri = icb_wcmd_attri_tmp;
  wire [1:0] icb_wcmd_xburst_tmp;
  assign icb_wcmd_xburst_tmp = wcmd_burst_r ? axi_awburst_buf : axi_awburst;
  assign icb_wcmd_xburst = icb_wcmd_xburst_tmp;
  wire [7:0] icb_wcmd_xlen_tmp;
  assign icb_wcmd_xlen_tmp = icb_wcmd_xburst_fixed ? 8'd0 : icb_wcmd_awlen;
  assign icb_wcmd_xlen = icb_wcmd_xlen_tmp;
  generate 
      if(ALLOW_FIX_BURST == 1) begin: allow_fix_burst_gen
  assign icb_wcmd_xburst_fixed = 1'b0;
      end
      else begin: disallow_fix_burst_gen
  assign icb_wcmd_xburst_fixed = (icb_wcmd_xburst == 2'b00);
      end
  endgenerate
endmodule
module  e603_subsys_gnrl_axi2ficb_r_id # (
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter USR_W = 4,
  parameter ID_W = 4
) (
  output                        icb_rrsp_ready,
  input                         icb_rrsp_valid,
  input [USR_W-1:0]             icb_rrsp_usr,
  input [DW-1:0]                icb_rrsp_rdata,
  input                         icb_rrsp_err,
  input                         icb_rrsp_excl_ok,
  input [ID_W-1:0]              icb_rrsp_id,
  input                         icb_rrsp_last,
  input                         axi_rready,
  output                        axi_rvalid,
  output [USR_W-1:0]            axi_ruser,
  output [ID_W-1:0]             axi_rid,
  output [DW-1:0]               axi_rdata,
  output [1:0]                  axi_rresp,
  output                        axi_rlast,
  input                         clk,
  input                         rst_n
  );
  assign icb_rrsp_ready   = axi_rready ;
  assign axi_rvalid       = icb_rrsp_valid ;
  wire [ID_W-1:0] axi_rid_tmp;
  assign axi_rid_tmp      = icb_rrsp_id;
  assign axi_rlast        = icb_rrsp_last;
  wire [DW-1:0] axi_rdata_tmp;
  assign axi_rdata_tmp    = icb_rrsp_rdata;
  assign axi_ruser        = icb_rrsp_usr;
  assign axi_rresp        = {icb_rrsp_err,icb_rrsp_excl_ok};
  assign axi_rdata = axi_rdata_tmp;
  assign axi_rid = axi_rid_tmp; 
endmodule
module  e603_subsys_gnrl_axi2ficb_b_id # (
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter USR_W = 4,
  parameter ID_W = 4
) (
  output                        icb_wrsp_ready,
  input                         icb_wrsp_valid,
  input                         icb_wrsp_err,
  input                         icb_wrsp_excl_ok,
  input [USR_W-1:0]             icb_wrsp_usr,
  input [ID_W-1:0]              icb_wrsp_id,
  input                         axi_bready,
  output                        axi_bvalid,
  output [1:0]                  axi_bresp,
  input [ID_W-1:0]             axi_bid,
  output [USR_W-1:0]             axi_buser,
  input [7:0]                   wrsp_xlen,
  input                         wrsp_burst,
  input                         wrsp_xlen_vld,
  input                         clk,
  input                         rst_n
  );
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_r_nxt;
  wire       burst_cnt_ena;
  assign burst_cnt_r_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_last = (burst_cnt_r == wrsp_xlen);
  assign burst_cnt_ena = wrsp_burst && icb_wrsp_valid && icb_wrsp_ready;
  assign icb_wrsp_ready   = ((wrsp_burst && !burst_last) || (axi_bready)) & wrsp_xlen_vld;
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_r_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign axi_bvalid = (icb_wrsp_valid && (!wrsp_burst || (wrsp_burst && burst_last))) & wrsp_xlen_vld;
  wire [1:0]  axi_bresp_nxt;
  wire [1:0]  axi_bresp_buf;
  wire        axi_bresp_en;
  assign axi_bresp_en = wrsp_burst && icb_wrsp_valid && icb_wrsp_ready && !burst_last;
  assign axi_bresp_nxt = (burst_cnt_r == 0) ? {icb_wrsp_err,icb_wrsp_excl_ok}
                                             : (axi_bresp_buf | {icb_wrsp_err,icb_wrsp_excl_ok})
                                             ;
e603_subsys_gnrl_dfflr #(2) bresp_dfflr (axi_bresp_en, axi_bresp_nxt, axi_bresp_buf, clk, rst_n);// VPP_NO_REG_PARSE
  assign axi_bresp = ({2{wrsp_burst}} & axi_bresp_buf) | {icb_wrsp_err,icb_wrsp_excl_ok};
  assign axi_buser = icb_wrsp_usr;
endmodule
module  e603_subsys_gnrl_axi2ficb_read_async_id # (
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 0,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input                            reset_flag_r,
  output                           axi_arready,
  input                            axi_arvalid,
  input [ID_W-1:0]                 axi_arid,
  input [AW-1:0]                   axi_araddr,
  input [7:0]                      axi_arlen,
  input [CMD_SIZE_W-1:0]                      axi_arsize,
  input [1:0]                      axi_arburst,
  input                            axi_arlock,
  input [3:0]                      axi_arcache,
  input [2:0]                      axi_arprot,
  input [USR_W-1:0]                axi_aruser,
  input                            axi_rready,
  output                           axi_rvalid,
  output [ID_W-1:0]                axi_rid,
  output [USR_W-1:0]               axi_ruser,
  output [DW-1:0]                  axi_rdata,
  output [1:0]                     axi_rresp,
  output                           axi_rlast,
  output                           icb_rcmd_sel   ,
  output                           icb_rcmd_valid ,
  input                            icb_rcmd_ready ,
  output [AW-1:0]                  icb_rcmd_addr  ,
  output                           icb_rcmd_read  ,
  output [DW-1:0]                  icb_rcmd_wdata ,
  output [MW-1:0]                  icb_rcmd_wmask ,
  output [1:0]                     icb_rcmd_beat  ,
  output                           icb_rcmd_excl  ,             
  output [CMD_SIZE_W-1:0]         icb_rcmd_size  ,
  output [7:0]                     icb_rcmd_xlen,
  output [1:0]                     icb_rcmd_xburst,
  output [1:0]                     icb_rcmd_modes,
  output                           icb_rcmd_dmode,
  output [2:0]                     icb_rcmd_attri,
  output [USR_W-1:0]               icb_rcmd_usr   ,
  output [ID_W-1:0]                icb_rcmd_id   ,
  output                           icb_rrsp_ready  , 
  input                            icb_rrsp_valid  , 
  input [DW-1:0]                   icb_rrsp_rdata  , 
  input [USR_W-1:0]                icb_rrsp_usr  , 
  input                            icb_rrsp_err    , 
  input                            icb_rrsp_excl_ok, 
  input [ID_W-1:0]                 icb_rrsp_id   ,
  input                            icb_rrsp_last,
  output                           axi2icb_read_axi_active,
  output                           axi2icb_read_icb_active,
  input icb_clk  ,
  input icb_rst_n,  
  input async_axi_clk  ,
  input async_axi_rst_n  
  );
  wire                           o_axi_arready;
  wire                           o_axi_arvalid;
  wire[ID_W-1:0]                 o_axi_arid;
  wire[AW-1:0]                   o_axi_araddr;
  wire[7:0]                      o_axi_arlen;
  wire[CMD_SIZE_W-1:0]                      o_axi_arsize;
  wire[1:0]                      o_axi_arburst;
  wire                           o_axi_arlock;
  wire[3:0]                      o_axi_arcache;
  wire[2:0]                      o_axi_arprot;
  wire[USR_W-1:0]                o_axi_aruser;
  wire                           o_axi_rready;
  wire                           o_axi_rvalid;
  wire [ID_W-1:0]                o_axi_rid;
  wire [USR_W-1:0]                o_axi_ruser;
  wire [DW-1:0]                  o_axi_rdata;
  wire [1:0]                     o_axi_rresp;
  wire                           o_axi_rlast;
  wire axi_buf_pipe_i_active;
  wire axi_buf_pipe_o_active;
  e603_subsys_gnrl_axi_buf_read # (
     .ASYNC (1),
     .SYNC_DP (SYNC_DP),
     .ASYNC_FIFO (ASYNC_FIFO),
     .ASYNC_FIFO_DP (ASYNC_FIFO_DP),
     .ASYNC_FIFO_DP_PTR_W (ASYNC_FIFO_DP_PTR_W),
     .RATIO_FIFO_DP(0),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW   (AW   ),
    .DW   (DW   ),
    .MW   (MW   ),
    .ID_W (ID_W ),
    .USR_W(USR_W) 
  ) u_axi_async_read(
    .reset_flag_r(reset_flag_r),
    .i_axi_arready        (axi_arready),
    .i_axi_arvalid        (axi_arvalid),
    .i_axi_arid           (axi_arid   ),
    .i_axi_araddr         (axi_araddr ),
    .i_axi_arlen          (axi_arlen  ),
    .i_axi_arsize         (axi_arsize ),
    .i_axi_arburst        (axi_arburst),
    .i_axi_arlock         (axi_arlock ),
    .i_axi_arcache        (axi_arcache),
    .i_axi_arprot         (axi_arprot ),
    .i_axi_aruser         (axi_aruser ),
    .i_axi_rready         (axi_rready ),
    .i_axi_rvalid         (axi_rvalid ),
    .i_axi_rid            (axi_rid    ),
    .i_axi_ruser          (axi_ruser    ),
    .i_axi_rdata          (axi_rdata  ),
    .i_axi_rresp          (axi_rresp  ),
    .i_axi_rlast          (axi_rlast  ),
    .o_axi_arready        (o_axi_arready),
    .o_axi_arvalid        (o_axi_arvalid),
    .o_axi_arid           (o_axi_arid   ),
    .o_axi_araddr         (o_axi_araddr ),
    .o_axi_arlen          (o_axi_arlen  ),
    .o_axi_arsize         (o_axi_arsize ),
    .o_axi_arburst        (o_axi_arburst),
    .o_axi_arlock         (o_axi_arlock ),
    .o_axi_arcache        (o_axi_arcache),
    .o_axi_arprot         (o_axi_arprot ),
    .o_axi_aruser         (o_axi_aruser ),
    .o_axi_rready         (o_axi_rready ),
    .o_axi_rvalid         (o_axi_rvalid ),
    .o_axi_rid            (o_axi_rid    ),
    .o_axi_ruser          (o_axi_ruser),
    .o_axi_rdata          (o_axi_rdata  ),
    .o_axi_rresp          (o_axi_rresp  ),
    .o_axi_rlast          (o_axi_rlast  ),
    .axi_buf_pipe_i_active  (axi_buf_pipe_i_active),
    .axi_buf_pipe_o_active  (axi_buf_pipe_o_active),
    .i_clk                (async_axi_clk  ),
    .i_rst_n              (async_axi_rst_n),
    .o_clk                (icb_clk  ),
    .o_rst_n              (icb_rst_n),
    .axi_bus_clk_en       (1'b1),
    .icb_clk_en           (1'b1),
    .clk                  (1'b0),
    .rst_n                (1'b0)  
  );
  wire o_axi2icb_read_active;
  e603_subsys_gnrl_axi2ficb_read_id # (
     .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
     .AW(AW),
     .DW(DW),
     .MW(MW),
     .RATIO_FIFO_DP(0),
     .FIFO_OUTS_NUM(FIFO_OUTS_NUM),
     .ID_W (ID_W),
     .USR_W (USR_W)
  ) u_axi2icb_read (
    .reset_flag_r    (1'b0),
    .axi_arready     (o_axi_arready ),
    .axi_arvalid     (o_axi_arvalid ),
    .axi_arid        (o_axi_arid    ),
    .axi_araddr      (o_axi_araddr  ),
    .axi_arlen       (o_axi_arlen   ),
    .axi_arsize      (o_axi_arsize  ),
    .axi_arburst     (o_axi_arburst ),
    .axi_arlock      (o_axi_arlock  ),
    .axi_arcache     (o_axi_arcache ),
    .axi_arprot      (o_axi_arprot  ),
    .axi_aruser      (o_axi_aruser  ),
    .axi_rready      (o_axi_rready   ),
    .axi_rvalid      (o_axi_rvalid   ),
    .axi_ruser       (o_axi_ruser    ),
    .axi_rid         (o_axi_rid      ),
    .axi_rdata       (o_axi_rdata    ),
    .axi_rresp       (o_axi_rresp    ),
    .axi_rlast       (o_axi_rlast    ),
    .icb_rcmd_sel    (icb_rcmd_sel    ),
    .icb_rcmd_valid  (icb_rcmd_valid  ),
    .icb_rcmd_ready  (icb_rcmd_ready  ),
    .icb_rcmd_addr   (icb_rcmd_addr   ),
    .icb_rcmd_read   (icb_rcmd_read   ),
    .icb_rcmd_wdata  (icb_rcmd_wdata  ),
    .icb_rcmd_wmask  (icb_rcmd_wmask  ),
    .icb_rcmd_beat   (icb_rcmd_beat   ),
    .icb_rcmd_excl   (icb_rcmd_excl   ),             
    .icb_rcmd_size   (icb_rcmd_size   ),
    .icb_rcmd_xlen   (icb_rcmd_xlen   ),
    .icb_rcmd_xburst (icb_rcmd_xburst ),
    .icb_rcmd_modes  (icb_rcmd_modes  ),
    .icb_rcmd_dmode  (icb_rcmd_dmode  ),
    .icb_rcmd_attri  (icb_rcmd_attri  ),
    .icb_rcmd_usr    (icb_rcmd_usr    ),
    .icb_rcmd_id     (icb_rcmd_id     ),
    .icb_rrsp_ready  (icb_rrsp_ready  ), 
    .icb_rrsp_valid  (icb_rrsp_valid  ), 
    .icb_rrsp_rdata  (icb_rrsp_rdata  ), 
    .icb_rrsp_err    (icb_rrsp_err    ), 
    .icb_rrsp_excl_ok(icb_rrsp_excl_ok), 
    .icb_rrsp_usr     (icb_rrsp_usr), 
    .icb_rrsp_id     (icb_rrsp_id), 
    .icb_rrsp_last   (icb_rrsp_last), 
    .axi_bus_clk_en  (1'b1),
    .icb_clk_en      (1'b1),
    .axi2icb_read_active  (o_axi2icb_read_active),
    .clk  (icb_clk  ),
    .rst_n(icb_rst_n)  
  );
  assign axi2icb_read_axi_active = axi_buf_pipe_i_active;
  assign axi2icb_read_icb_active = axi_buf_pipe_o_active | o_axi2icb_read_active;
endmodule
module  e603_subsys_gnrl_axi2ficb_write_async_id # (
  parameter ALLOW_FIX_BURST = 0,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 0,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           axi_awready,
  input                            axi_awvalid,
  input [ID_W-1:0]                 axi_awid,
  input [AW-1:0]                   axi_awaddr,
  input [7:0]                      axi_awlen,
  input [CMD_SIZE_W-1:0]                      axi_awsize,
  input [1:0]                      axi_awburst,
  input                            axi_awlock,
  input [3:0]                      axi_awcache,
  input [2:0]                      axi_awprot,
  input [USR_W-1:0]                axi_awuser, 
  output                           axi_wready,
  input                            axi_wvalid,
  input [DW-1:0]                   axi_wdata,
  input [MW-1:0]                   axi_wstrb,
  input                            axi_wlast,
  input                            axi_bready,
  output                           axi_bvalid,
  output [USR_W-1:0]               axi_buser,
  output [ID_W-1:0]                axi_bid,
  output [1:0]                     axi_bresp,
  output                           icb_wcmd_sel,
  output                           icb_wcmd_valid,
  input                            icb_wcmd_ready,
  output [AW-1:0]                  icb_wcmd_addr,
  output                           icb_wcmd_read, 
  output [DW-1:0]                  icb_wcmd_wdata,
  output [MW-1:0]                  icb_wcmd_wmask,
  output [1:0]                     icb_wcmd_beat,
  output                           icb_wcmd_lock,
  output                           icb_wcmd_excl,
  output [CMD_SIZE_W-1:0]         icb_wcmd_size,
  output [7:0]                     icb_wcmd_xlen,
  output [1:0]                     icb_wcmd_xburst,
  output [1:0]                     icb_wcmd_modes,
  output                           icb_wcmd_dmode,
  output [2:0]                     icb_wcmd_attri,
  output [USR_W-1:0]               icb_wcmd_usr,
  output [ID_W-1:0]                icb_wcmd_id,
  input                            icb_wrsp_valid,
  output                           icb_wrsp_ready,
  input                            icb_wrsp_err,
  input                            icb_wrsp_excl_ok,
  input [USR_W-1:0]                icb_wrsp_usr,
  input [ID_W-1:0]                 icb_wrsp_id,
  output                           axi2icb_write_axi_active,
  output                           axi2icb_write_icb_active,
  input icb_clk  ,
  input icb_rst_n,  
  input async_axi_clk  ,
  input async_axi_rst_n  
  );
  wire                           o_axi_awready;
  wire                           o_axi_awvalid;
  wire[ID_W-1:0]                 o_axi_awid;
  wire[AW-1:0]                   o_axi_awaddr;
  wire[7:0]                      o_axi_awlen;
  wire[CMD_SIZE_W-1:0]                      o_axi_awsize;
  wire[1:0]                      o_axi_awburst;
  wire                           o_axi_awlock;
  wire[3:0]                      o_axi_awcache;
  wire[2:0]                      o_axi_awprot;
  wire[USR_W-1:0]                o_axi_awuser; 
  wire                           o_axi_wready;
  wire                           o_axi_wvalid;
  wire[DW-1:0]                   o_axi_wdata;
  wire[MW-1:0]                   o_axi_wstrb;
  wire                           o_axi_wlast;
  wire                           o_axi_bready;
  wire                           o_axi_bvalid;
  wire [USR_W-1:0]               o_axi_buser;
  wire [ID_W-1:0]                o_axi_bid;
  wire [1:0]                     o_axi_bresp;
  wire axi_buf_pipe_i_active;
  wire axi_buf_pipe_o_active;
  e603_subsys_gnrl_axi_buf_write # (
     .ASYNC (1),
     .SYNC_DP (SYNC_DP),
     .ASYNC_FIFO (ASYNC_FIFO),
     .ASYNC_FIFO_DP (ASYNC_FIFO_DP),
     .ASYNC_FIFO_DP_PTR_W (ASYNC_FIFO_DP_PTR_W),
     .RATIO_FIFO_DP(0),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW   (AW   ),
    .DW   (DW   ),
    .MW   (MW   ),
    .ID_W (ID_W ),
    .USR_W(USR_W) 
  ) u_axi_buf_write (
    .reset_flag_r(reset_flag_r),
    .i_axi_awready   (axi_awready   ),
    .i_axi_awvalid   (axi_awvalid   ),
    .i_axi_awid      (axi_awid      ),
    .i_axi_awaddr    (axi_awaddr    ),
    .i_axi_awlen     (axi_awlen     ),
    .i_axi_awsize    (axi_awsize    ),
    .i_axi_awburst   (axi_awburst   ),
    .i_axi_awlock    (axi_awlock    ),
    .i_axi_awcache   (axi_awcache   ),
    .i_axi_awprot    (axi_awprot    ),
    .i_axi_awuser    (axi_awuser    ), 
    .i_axi_wready    (axi_wready    ),
    .i_axi_wvalid    (axi_wvalid    ),
    .i_axi_wdata     (axi_wdata     ),
    .i_axi_wstrb     (axi_wstrb     ),
    .i_axi_wlast     (axi_wlast     ),
    .i_axi_bready    (axi_bready    ),
    .i_axi_bvalid    (axi_bvalid    ),
    .i_axi_buser     (axi_buser     ),
    .i_axi_bid       (axi_bid       ),
    .i_axi_bresp     (axi_bresp     ),
    .o_axi_awready   (o_axi_awready   ),
    .o_axi_awvalid   (o_axi_awvalid   ),
    .o_axi_awid      (o_axi_awid      ),
    .o_axi_awaddr    (o_axi_awaddr    ),
    .o_axi_awlen     (o_axi_awlen     ),
    .o_axi_awsize    (o_axi_awsize    ),
    .o_axi_awburst   (o_axi_awburst   ),
    .o_axi_awlock    (o_axi_awlock    ),
    .o_axi_awcache   (o_axi_awcache   ),
    .o_axi_awprot    (o_axi_awprot    ),
    .o_axi_awuser    (o_axi_awuser    ), 
    .o_axi_wready    (o_axi_wready    ),
    .o_axi_wvalid    (o_axi_wvalid    ),
    .o_axi_wdata     (o_axi_wdata     ),
    .o_axi_wstrb     (o_axi_wstrb     ),
    .o_axi_wlast     (o_axi_wlast     ),
    .o_axi_bready    (o_axi_bready    ),
    .o_axi_bvalid    (o_axi_bvalid    ),
    .o_axi_bid       (o_axi_bid       ),
    .o_axi_buser     (o_axi_buser     ),
    .o_axi_bresp     (o_axi_bresp     ),
    .axi_buf_pipe_i_active  (axi_buf_pipe_i_active),
    .axi_buf_pipe_o_active  (axi_buf_pipe_o_active),
    .i_clk                (async_axi_clk  ),
    .i_rst_n              (async_axi_rst_n),
    .o_clk                (icb_clk  ),
    .o_rst_n              (icb_rst_n),
    .axi_bus_clk_en       (1'b1),
    .icb_clk_en       (1'b1),
    .clk                  (1'b0),
    .rst_n                (1'b0)  
  );
  wire o_axi2icb_write_active;
  e603_subsys_gnrl_axi2ficb_write_id # (
  .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
  .AW(AW),
  .DW(DW),
  .MW(MW),
  .RATIO_FIFO_DP(0),
  .FIFO_OUTS_NUM(FIFO_OUTS_NUM),
  .ID_W (ID_W),
  .USR_W (USR_W)
  ) u_axi2icb_write (
    .reset_flag_r (1'b0),
    .axi_awready   (o_axi_awready   ),
    .axi_awvalid   (o_axi_awvalid   ),
    .axi_awid      (o_axi_awid      ),
    .axi_awaddr    (o_axi_awaddr    ),
    .axi_awlen     (o_axi_awlen     ),
    .axi_awsize    (o_axi_awsize    ),
    .axi_awburst   (o_axi_awburst   ),
    .axi_awlock    (o_axi_awlock    ),
    .axi_awcache   (o_axi_awcache   ),
    .axi_awprot    (o_axi_awprot    ),
    .axi_awuser    (o_axi_awuser    ), 
    .axi_wready    (o_axi_wready    ),
    .axi_wvalid    (o_axi_wvalid    ),
    .axi_wdata     (o_axi_wdata     ),
    .axi_wstrb     (o_axi_wstrb     ),
    .axi_wlast     (o_axi_wlast     ),
    .axi_bready    (o_axi_bready    ),
    .axi_bvalid    (o_axi_bvalid    ),
    .axi_bid       (o_axi_bid       ),
    .axi_buser     (o_axi_buser     ),
    .axi_bresp     (o_axi_bresp     ),
    .icb_wcmd_sel   (icb_wcmd_sel),
    .icb_wcmd_valid (icb_wcmd_valid ),
    .icb_wcmd_ready (icb_wcmd_ready ),
    .icb_wcmd_addr  (icb_wcmd_addr  ),
    .icb_wcmd_read  (icb_wcmd_read  ), 
    .icb_wcmd_wdata (icb_wcmd_wdata ),
    .icb_wcmd_wmask (icb_wcmd_wmask ),
    .icb_wcmd_beat  (icb_wcmd_beat  ),
    .icb_wcmd_lock  (icb_wcmd_lock  ),
    .icb_wcmd_excl  (icb_wcmd_excl  ),
    .icb_wcmd_size  (icb_wcmd_size  ),
    .icb_wcmd_xlen  (icb_wcmd_xlen    ),
    .icb_wcmd_xburst(icb_wcmd_xburst  ),
    .icb_wcmd_modes (icb_wcmd_modes   ),
    .icb_wcmd_dmode (icb_wcmd_dmode   ),
    .icb_wcmd_attri (icb_wcmd_attri   ),
    .icb_wcmd_usr   (icb_wcmd_usr ),
    .icb_wcmd_id    (icb_wcmd_id),
    .icb_wrsp_valid  (icb_wrsp_valid  ),
    .icb_wrsp_ready  (icb_wrsp_ready  ),
    .icb_wrsp_err    (icb_wrsp_err    ),
    .icb_wrsp_excl_ok(icb_wrsp_excl_ok),
    .icb_wrsp_id     (icb_wrsp_id),
    .icb_wrsp_usr     (icb_wrsp_usr),
    .axi_bus_clk_en  (1'b1),
    .icb_clk_en  (1'b1),
    .axi2icb_write_active  (o_axi2icb_write_active),
    .clk   (icb_clk  ),
    .rst_n (icb_rst_n)
  );
  assign axi2icb_write_axi_active = axi_buf_pipe_i_active;
  assign axi2icb_write_icb_active = axi_buf_pipe_o_active | o_axi2icb_write_active;
endmodule
`include "global.v"
module e603_subsys_gnrl_ficb2axi_ar # (
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_UW = 1 
) (
  output                        ar_pend_active,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input                         icb_cmd_read, 
  input [AW-1:0]                icb_cmd_addr, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input                         axi_arready,
  output                        axi_arvalid,
  output [AW-1:0]               axi_araddr,
  output [AXLEN_W-1:0]                  axi_arlen,
  output [CMD_SIZE_W-1:0]                  axi_arsize,
  output [1:0]                  axi_arburst,
  output                        axi_arlock,
  output [3:0]                  axi_arcache,
  output [2:0]                  axi_arprot,
  output [CMD_UW-1:0]            axi_aruser,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_W = AW+AXLEN_W+CMD_SIZE_W+1+2+4+3+CMD_UW 
                    ;
  wire              i_arvalid;
  wire [AW-1:0]     i_araddr;
  wire [AXLEN_W-1:0]        i_arlen;
  wire [CMD_SIZE_W-1:0]        i_arsize;
  wire [1:0]        i_arburst;
  wire              i_arlock;
  wire [3:0]        i_arcache;
  wire [2:0]        i_arprot;
  wire [CMD_UW-1:0]  i_aruser;
  wire [PACK_W-1:0] i_axi_pack;
  wire [PACK_W-1:0] o_axi_pack;
  wire i_axi_vld;
  wire i_axi_rdy;
  wire o_axi_vld;
  wire o_axi_rdy;
  wire axi_ar_ready;
  wire burst_flag_r;
  wire burst_flag_en;
  wire burst_flag_set;
  wire burst_flag_clr;
  assign burst_flag_en = burst_flag_set || burst_flag_clr;
  assign axi_ar_ready = axi_arready;
  assign burst_flag_set = icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[0] & icb_clk_en;
  assign burst_flag_clr = burst_flag_r && icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[1] & icb_clk_en;
e603_subsys_gnrl_dfflr #(1) burst_flag_dfflr (burst_flag_en, burst_flag_set, burst_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign ar_pend_active = burst_flag_r;
  assign icb_cmd_ready = i_axi_rdy | burst_flag_r;
  assign i_arvalid = icb_cmd_valid & (~burst_flag_r);
  assign i_araddr   = icb_cmd_addr;
  assign i_arlen     = icb_cmd_xlen[AXLEN_W-1:0];
  assign i_arburst   = ((icb_cmd_xlen == {AXLEN_W{1'b0}}) & (icb_cmd_xburst[1:0] == 2'b0)) ? 2'b01 : icb_cmd_xburst[1:0];
  assign i_arsize    = icb_cmd_size;
  assign i_arlock    = icb_cmd_excl; 
  wire icb_cmd_mmode  = (icb_cmd_modes == 2'd0);
  wire icb_cmd_smode  = (icb_cmd_modes == 2'd2);
  wire icb_cmd_ifu    = icb_cmd_attri[0];
  wire icb_cmd_device = icb_cmd_attri[1];
  wire icb_cmd_nc     = icb_cmd_attri[2];
  assign i_arcache   =  (icb_cmd_device & icb_cmd_nc) ? 4'b1011 : 
                        icb_cmd_device ? 4'b0000 :
                        icb_cmd_nc     ? 4'b0011 : 4'b1111;
  assign i_arprot[0] = icb_cmd_mmode;
  assign i_arprot[1] = 1'b0; 
  assign i_arprot[2] = icb_cmd_ifu;
  assign i_aruser    = icb_cmd_usr;
  assign i_axi_pack = 
                      {
                        i_araddr,
                        i_arlen,
                        i_arsize,
                        i_arburst,
                        i_arlock,
                        i_arcache,
                        i_arprot,
                        i_aruser 
                      };
  assign {
           axi_araddr,
           axi_arlen,
           axi_arsize,
           axi_arburst,
           axi_arlock,
           axi_arcache,
           axi_arprot,
           axi_aruser 
         } = o_axi_pack;
  assign axi_arvalid = o_axi_vld;
  assign i_axi_vld = i_arvalid;
  assign o_axi_rdy = axi_ar_ready;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_W)
  ) u_axi_ar_fifo (
        .i_clk_en(icb_clk_en),
        .i_vld(i_axi_vld),
        .i_rdy(i_axi_rdy),
        .i_dat(i_axi_pack),
        .o_clk_en(axi_bus_clk_en),
        .o_vld(o_axi_vld),
        .o_rdy(o_axi_rdy),  
        .o_dat(o_axi_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb2axi_aw # (
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_UW = 1
) (
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input                         axi_awready,
  output                        axi_awvalid,
  output [AW-1:0]               axi_awaddr,
  output [AXLEN_W-1:0]                  axi_awlen,
  output [CMD_SIZE_W-1:0]                  axi_awsize,
  output [1:0]                  axi_awburst,
  output                        axi_awlock,
  output [3:0]                  axi_awcache,
  output [2:0]                  axi_awprot,
  output [CMD_UW-1:0]            axi_awuser, 
  input                         axi_wready,
  output                        axi_wvalid,
  output [DW-1:0]               axi_wdata,
  output [DW/8-1:0]               axi_wstrb,
  output                        axi_wlast,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_A_W = AW+AXLEN_W+CMD_SIZE_W+1+2+4+3+CMD_UW 
                           ;
  localparam PACK_D_W = DW+DW/8+1;
  wire axi_aw_ready;
  wire axi_w_ready;
  wire burst_flag_r;
  wire burst_flag_en;
  wire burst_flag_set;
  wire burst_flag_clr;
  wire [PACK_A_W-1:0] i_axi_a_pack;
  wire [PACK_A_W-1:0] o_axi_a_pack;
  wire [PACK_D_W-1:0] i_axi_d_pack;
  wire [PACK_D_W-1:0] o_axi_d_pack;
  wire i_axi_a_vld;
  wire i_axi_a_rdy;
  wire o_axi_a_vld;
  wire o_axi_a_rdy;
  wire i_axi_d_vld;
  wire i_axi_d_rdy;
  wire o_axi_d_vld;
  wire o_axi_d_rdy;
  wire                i_awready;
  wire                i_awvalid;
  wire [AW-1:0]       i_awaddr;
  wire [AXLEN_W-1:0]          i_awlen;
  wire [CMD_SIZE_W-1:0]          i_awsize;
  wire [1:0]          i_awburst;
  wire                i_awlock;
  wire [3:0]          i_awcache;
  wire [2:0]          i_awprot;
  wire [CMD_UW-1:0]    i_awuser; 
  wire                i_wready;
  wire                i_wvalid;
  wire [DW-1:0]       i_wdata;
  wire [DW/8-1:0]       i_wstrb;
  wire                i_wlast;
  assign axi_aw_ready = axi_awready ;
  assign axi_w_ready  = axi_wready  ;
  assign i_axi_a_pack = 
                      {
                        i_awaddr,
                        i_awlen,
                        i_awsize,
                        i_awburst,
                        i_awlock,
                        i_awcache,
                        i_awprot,
                        i_awuser  
                      };
  assign i_axi_a_vld = i_awvalid;
  assign i_awready = i_axi_a_rdy; 
  assign {
          axi_awaddr,
          axi_awlen,
          axi_awsize,
          axi_awburst,
          axi_awlock,
          axi_awcache,
          axi_awprot,
          axi_awuser  
         } = o_axi_a_pack;
  assign axi_awvalid = o_axi_a_vld;
  assign o_axi_a_rdy = axi_aw_ready;
  assign i_axi_d_pack = 
                      {
                       i_wdata,
                       i_wstrb,
                       i_wlast
                      };
  assign i_axi_d_vld = i_wvalid;
  assign i_wready    = i_axi_d_rdy; 
  assign {
          axi_wdata,
          axi_wstrb,
          axi_wlast
         } = o_axi_d_pack;
  assign axi_wvalid  = o_axi_d_vld;
  assign o_axi_d_rdy = axi_w_ready;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_A_W)
  ) u_axi_aw_fifo (
        .i_clk_en(icb_clk_en),
        .i_vld(i_axi_a_vld),
        .i_rdy(i_axi_a_rdy),
        .i_dat(i_axi_a_pack),
        .o_clk_en(axi_bus_clk_en),
        .o_vld(o_axi_a_vld),
        .o_rdy(o_axi_a_rdy),  
        .o_dat(o_axi_a_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_D_W)
  ) u_axi_w_fifo (
        .i_clk_en(icb_clk_en),
        .i_vld(i_axi_d_vld),
        .i_rdy(i_axi_d_rdy),
        .i_dat(i_axi_d_pack),
        .o_clk_en(axi_bus_clk_en),
        .o_vld(o_axi_d_vld),
        .o_rdy(o_axi_d_rdy),  
        .o_dat(o_axi_d_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  assign burst_flag_en = burst_flag_set || burst_flag_clr;
  assign burst_flag_set = icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[0] & icb_clk_en
                        ;
  assign burst_flag_clr = burst_flag_r && icb_cmd_ready && icb_cmd_valid && icb_cmd_beat[1] & icb_clk_en;
e603_subsys_gnrl_dfflr #(1) burst_flag_dfflr (burst_flag_en, burst_flag_set, burst_flag_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_cmd_ready =   (i_awready || burst_flag_r) && (i_wready);
  assign i_awvalid = icb_cmd_valid && (!burst_flag_r) && i_wready;
  assign i_wvalid  = icb_cmd_valid && (i_awready || burst_flag_r);
  assign i_awaddr   = icb_cmd_addr;
  assign i_awlen     = icb_cmd_xlen[AXLEN_W-1:0];
  assign i_awburst   = ((icb_cmd_xlen == {AXLEN_W{1'b0}}) & (icb_cmd_xburst[1:0] == 2'b0)) ? 2'b01 : icb_cmd_xburst[1:0];
  assign i_awsize    = icb_cmd_size;
  assign i_awlock    = icb_cmd_excl; 
  wire icb_cmd_mmode  = (icb_cmd_modes == 2'd0);
  wire icb_cmd_smode  = (icb_cmd_modes == 2'd2);
  wire icb_cmd_ifu    = icb_cmd_attri[0];
  wire icb_cmd_device = icb_cmd_attri[1];
  wire icb_cmd_nc     = icb_cmd_attri[2];
  assign i_awcache   =  (icb_cmd_device & icb_cmd_nc) ? 4'b0111 : 
                        icb_cmd_device ? 4'b0000 :
                          icb_cmd_nc     ? 4'b0011 : 4'b1111;
  assign i_awprot[0] = icb_cmd_mmode;
  assign i_awprot[1] = 1'b0; 
  assign i_awprot[2] = 1'b0;
  assign i_awuser    = icb_cmd_usr;
  assign i_wdata     = icb_cmd_wdata;
  assign i_wstrb     = icb_cmd_wmask;   
  assign i_wlast    = ((icb_cmd_beat == 2'b00) && !burst_flag_r) || icb_cmd_beat[1];
endmodule
module e603_subsys_gnrl_ficb2axi_r # (
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter REG_OUT = 0,
  parameter RSP_UW = 1 
) (
  input                          icb_cmd_cnt_is_0,
  output                         icb_rrsp_valid,
  input                          icb_rrsp_ready,
  output [DW-1:0]                icb_rrsp_rdata,
  output                         icb_rrsp_err,
  output                         icb_rrsp_excl_ok,
  output [RSP_UW-1:0]            icb_rrsp_usr,
  output                         axi_rready,
  input                          axi_rvalid,
  input [RSP_UW-1:0]              axi_ruser,
  input [DW-1:0]                 axi_rdata,
  input [1:0]                    axi_rresp,
  input                          axi_rlast,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_W = DW+2+1+RSP_UW;
  wire                          o_rvalid;
  wire [DW-1:0]                 o_rdata;
  wire [RSP_UW-1:0]              o_rusr;
  wire [1:0]                    o_rresp;
  wire                          o_rlast;
  wire [PACK_W-1:0] i_axi_pack;
  wire [PACK_W-1:0] o_axi_pack;
  wire i_axi_vld;
  wire i_axi_rdy;
  wire o_axi_vld;
  wire o_axi_rdy;
  assign i_axi_pack = 
                      {
                        axi_ruser,
                        axi_rdata,
                        axi_rresp,
                        axi_rlast 
                      };
  assign {
          o_rusr,
          o_rdata,
          o_rresp,
          o_rlast 
         } = o_axi_pack;
  assign o_rvalid = o_axi_vld;
  assign icb_rrsp_valid = (~icb_cmd_cnt_is_0) & o_rvalid      ;
  assign o_axi_rdy      = (~icb_cmd_cnt_is_0) & icb_rrsp_ready;
  assign i_axi_vld = axi_rvalid ;
  assign axi_rready = i_axi_rdy;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .REG_OUT (REG_OUT),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_W)
  ) u_axi_r_fifo (
        .i_clk_en(axi_bus_clk_en),
        .i_vld(i_axi_vld),
        .i_rdy(i_axi_rdy),
        .i_dat(i_axi_pack),
        .o_clk_en(icb_clk_en),
        .o_vld(o_axi_vld),
        .o_rdy(o_axi_rdy),  
        .o_dat(o_axi_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  wire icb_rrsp_err_tmp     = o_rresp[1]   
                 ;
  assign icb_rrsp_err = icb_rrsp_err_tmp;
  wire icb_rrsp_excl_ok_tmp = (o_rresp == 2'b01);
  assign icb_rrsp_excl_ok = icb_rrsp_excl_ok_tmp;
  assign icb_rrsp_rdata   = o_rdata;
  assign icb_rrsp_usr     = o_rusr;
endmodule
module e603_subsys_gnrl_ficb2axi_b # (
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter RSP_UW = 1,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2 
) (
  input                          wrsp_burst_fifo_o_vld,
  output                         icb_wrsp_valid,
  input                          icb_wrsp_ready,
  output                         icb_wrsp_err,
  output                         icb_wrsp_excl_ok,
  output [RSP_UW-1:0]             icb_wrsp_usr,
  output                         axi_bready,
  input                          axi_bvalid,
  input [1:0]                    axi_bresp,
  input [RSP_UW-1:0]              axi_buser,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input [7:0]                   wrsp_xlen,
  output                        wrsp_last,
  input                         clk,
  input                         rst_n
  );
  localparam PACK_W = 2+RSP_UW;
  wire [RSP_UW-1:0]              o_busr;
  wire [1:0]                    o_bresp;
  wire o_burst = (wrsp_xlen != 8'b0);
  wire [PACK_W-1:0] i_axi_pack;
  wire [PACK_W-1:0] o_axi_pack;
  wire i_axi_vld;
  wire i_axi_rdy;
  wire o_axi_vld;
  wire o_axi_rdy;
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_r_nxt;
  wire       burst_cnt_ena;
  assign i_axi_pack = 
                      {
                        axi_bresp,
                        axi_buser 
                      };
  assign {
          o_bresp,
          o_busr 
         } = o_axi_pack;
  assign i_axi_vld = axi_bvalid ;
  assign axi_bready = i_axi_rdy;
  e603_subsys_gnrl_ratio_fifo # (
        .I_SUPPORT_RATIO (1),
        .O_SUPPORT_RATIO (1),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DP  (RATIO_FIFO_DP),
        .DW  (PACK_W)
  ) u_axi_b_fifo (
        .i_clk_en(axi_bus_clk_en),
        .i_vld(i_axi_vld),
        .i_rdy(i_axi_rdy),
        .i_dat(i_axi_pack),
        .o_clk_en(icb_clk_en),
        .o_vld(o_axi_vld),
        .o_rdy(o_axi_rdy),  
        .o_dat(o_axi_pack),  
        .o_fifo_active(),
        .clk  (clk),
        .rst_n(rst_n)
  );
  wire burst_first = (burst_cnt_r == 8'd0);
  assign burst_cnt_r_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_cnt_ena = o_burst && icb_wrsp_valid && icb_wrsp_ready & icb_clk_en;
  assign burst_last = (burst_cnt_r == wrsp_xlen) & (~burst_first);
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_r_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_wrsp_valid   = wrsp_last ? o_axi_vld : wrsp_burst_fifo_o_vld;
  assign o_axi_rdy = icb_wrsp_ready && wrsp_last;
  wire icb_wrsp_err_tmp     = wrsp_last ? (o_bresp[1] 
                                        ): 1'b0;
  assign icb_wrsp_err     = icb_wrsp_err_tmp;
  wire icb_wrsp_excl_ok_tmp = wrsp_last ? (o_bresp == 2'b01) : 1'b0;
  assign icb_wrsp_excl_ok = icb_wrsp_excl_ok_tmp;
  assign icb_wrsp_usr     = wrsp_last ? o_busr : {RSP_UW{1'b0}};
  assign wrsp_last = burst_last | (wrsp_xlen == 8'd0);
   endmodule
module e603_subsys_gnrl_ficb2axi_read # (
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter REG_OUT = 0,
  parameter OUTS_CNT_W = 4,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  output icb2axi_read_pend_active,
  input                         axi_arready,
  output                        axi_arvalid,
  output [AW-1:0]               axi_araddr,
  output [AXLEN_W-1:0]                  axi_arlen,
  output [CMD_SIZE_W-1:0]                  axi_arsize,
  output [1:0]                  axi_arburst,
  output                        axi_arlock,
  output [3:0]                  axi_arcache,
  output [2:0]                  axi_arprot,
  output [CMD_UW-1:0]            axi_aruser,
  output                        axi_rready,
  input                         axi_rvalid,
  input [DW-1:0]                axi_rdata,
  input [RSP_UW-1:0]             axi_ruser,
  input [1:0]                   axi_rresp,
  input                         axi_rlast,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]            icb_rsp_usr,
  input                         clk,
  input                         rst_n
  );
  localparam CNT_W = 8;
  wire outs_cnt_inc = icb_cmd_valid & icb_cmd_ready & icb_clk_en;
  wire outs_cnt_dec = icb_rsp_valid & icb_rsp_ready & icb_clk_en;
  wire outs_cnt_ena = outs_cnt_inc ^ outs_cnt_dec;
  wire [CNT_W-1:0] outs_cnt_r;
  wire [CNT_W-1:0] outs_cnt_nxt = outs_cnt_inc ? (outs_cnt_r + 1'b1) : (outs_cnt_r - 1'b1);
e603_subsys_gnrl_dfflr #(CNT_W) outs_cnt_dfflr (outs_cnt_ena, outs_cnt_nxt, outs_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  wire icb_cmd_cnt_full = (outs_cnt_r == {CNT_W{1'b1}});
  wire icb_cmd_cnt_is_0 = (outs_cnt_r == {CNT_W{1'b0}});
  wire icb_cmd_valid_raw;
  wire icb_cmd_ready_raw;
  assign icb_cmd_valid_raw = (~icb_cmd_cnt_full) & icb_cmd_valid;
  assign icb_cmd_ready     = (~icb_cmd_cnt_full) & icb_cmd_ready_raw;
  wire ar_pend_active;
  assign icb2axi_read_pend_active = (~icb_cmd_cnt_is_0) | ar_pend_active | axi_arvalid;
 e603_subsys_gnrl_ficb2axi_ar # (
            .AXLEN_W (AXLEN_W),
            .AW (AW),
            .DW (DW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP),
            .CMD_SIZE_W(CMD_SIZE_W),
            .CMD_UW (CMD_UW)
   ) u_icb2axi_ar(
            .ar_pend_active(ar_pend_active),
            .icb_cmd_valid (icb_cmd_valid_raw),
            .icb_cmd_ready (icb_cmd_ready_raw),
            .icb_cmd_addr (icb_cmd_addr), 
            .icb_cmd_sel  (icb_cmd_sel), 
            .icb_cmd_xlen(icb_cmd_xlen),
            .icb_cmd_xburst(icb_cmd_xburst),
            .icb_cmd_modes (icb_cmd_modes ),
            .icb_cmd_dmode (icb_cmd_dmode ),
            .icb_cmd_attri (icb_cmd_attri ),
            .icb_cmd_read (icb_cmd_read), 
            .icb_cmd_wdata (icb_cmd_wdata),
            .icb_cmd_wmask (icb_cmd_wmask),
            .icb_cmd_beat (icb_cmd_beat),
            .icb_cmd_lock (icb_cmd_lock),
            .icb_cmd_excl (icb_cmd_excl),
            .icb_cmd_size (icb_cmd_size),
            .icb_cmd_usr (icb_cmd_usr),
            .axi_arready (axi_arready),
            .axi_arvalid (axi_arvalid),
            .axi_araddr (axi_araddr),
            .axi_arlen (axi_arlen),
            .axi_arsize (axi_arsize),
            .axi_arburst (axi_arburst),
            .axi_arlock (axi_arlock),
            .axi_arcache (axi_arcache),
            .axi_arprot (axi_arprot),
            .axi_aruser (axi_aruser),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .clk (clk),
            .rst_n (rst_n)
  );
  e603_subsys_gnrl_ficb2axi_r # (
            .AW (AW),
            .DW (DW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP),
            .REG_OUT(REG_OUT),
            .RSP_UW (RSP_UW) 
  ) u_icb2axi_r(
            .icb_cmd_cnt_is_0(icb_cmd_cnt_is_0),
            .icb_rrsp_valid (icb_rsp_valid),
            .icb_rrsp_ready (icb_rsp_ready),
            .icb_rrsp_rdata (icb_rsp_rdata),
            .icb_rrsp_usr (icb_rsp_usr),
            .icb_rrsp_err (icb_rsp_err),
            .icb_rrsp_excl_ok (icb_rsp_excl_ok),
            .axi_rready (axi_rready),
            .axi_rvalid (axi_rvalid),
            .axi_rdata (axi_rdata),
            .axi_ruser (axi_ruser),
            .axi_rresp (axi_rresp),
            .axi_rlast (axi_rlast),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .clk (clk),
            .rst_n (rst_n)
  );
endmodule
module e603_subsys_gnrl_ficb2axi_write # (
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter OUTS_CNT_W =2,
  parameter SUPPORT_AWID_OOO = 0,
  parameter OUTS_FIFO_DP =4,
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP =2,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
) (
  output                        icb2axi_write_pend_active,
  input                         axi_awready,
  output                        axi_awvalid,
  output [AW-1:0]               axi_awaddr,
  output [AXLEN_W-1:0]                  axi_awlen,
  output [CMD_SIZE_W-1:0]                  axi_awsize,
  output [1:0]                  axi_awburst,
  output                        axi_awlock,
  output [3:0]                  axi_awcache,
  output [2:0]                  axi_awprot,
  output [CMD_UW-1:0]            axi_awuser, 
  input                         axi_wready,
  output                        axi_wvalid,
  output [DW-1:0]               axi_wdata,
  output [DW/8-1:0]               axi_wstrb,
  output                        axi_wlast,
  output                         axi_bready,
  input                          axi_bvalid,
  input [RSP_UW-1:0]              axi_buser,
  input [1:0]                    axi_bresp,
  input                         axi_bus_clk_en,
  input                         icb_clk_en,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr,
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [AXLEN_W-1:0]                   icb_cmd_xlen,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err,
  output                        icb_rsp_excl_ok,
  output[RSP_UW-1:0]             icb_rsp_usr,
  output[DW-1:0]                icb_rsp_rdata,
  input                         clk,
  input                         rst_n
  );
  assign icb_rsp_rdata = {DW{1'b0}};
  wire [7:0] wrsp_xlen;
  wire [7:0] wcmd_xlen;
  wire wrsp_burst_fifo_i_vld;
  wire wrsp_burst_fifo_o_rdy;
  wire wrsp_burst_fifo_o_vld;
  wire wrsp_burst_fifo_i_rdy;
  wire wrsp_last;
  wire icb_cmd_valid_raw;
  wire icb_cmd_ready_raw;
  assign icb_cmd_valid_raw = wrsp_burst_fifo_i_rdy & icb_cmd_valid;
  assign icb_cmd_ready     = wrsp_burst_fifo_i_rdy & icb_cmd_ready_raw;
  assign wrsp_burst_fifo_i_vld = icb_cmd_valid & icb_cmd_ready;
  assign wrsp_burst_fifo_o_rdy = icb_rsp_valid & icb_rsp_ready;
  assign wcmd_xlen = icb_cmd_xlen[7:0];
  generate
    if(SUPPORT_AWID_OOO == 1) begin: ooo_is1
  e603_subsys_gnrl_fifo # (
        .REG_OUT(1),
        .DP  (OUTS_FIFO_DP),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DW  (8)
  ) u_wrsp_burst_fifo (
        .i_vld(wrsp_burst_fifo_i_vld & icb_clk_en),
        .i_rdy(wrsp_burst_fifo_i_rdy),
        .i_dat(wcmd_xlen),
        .o_vld(wrsp_burst_fifo_o_vld),
        .o_rdy(wrsp_burst_fifo_o_rdy & icb_clk_en),  
        .o_dat(wrsp_xlen),  
        .clk  (clk),
        .rst_n(rst_n)
  );
    end
    else begin: ooo_is0
     e603_subsys_gnrl_fifo # (
        .REG_OUT(1),
        .DP  (OUTS_FIFO_DP),
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .DW  (8)
  ) u_wrsp_burst_fifo (
        .i_vld(wrsp_burst_fifo_i_vld & icb_clk_en),
        .i_rdy(wrsp_burst_fifo_i_rdy),
        .i_dat(wcmd_xlen),
        .o_vld(wrsp_burst_fifo_o_vld),
        .o_rdy(wrsp_burst_fifo_o_rdy & icb_clk_en),  
        .o_dat(wrsp_xlen),  
        .clk  (clk),
        .rst_n(rst_n)
  );
    end
  endgenerate
 e603_subsys_gnrl_ficb2axi_aw # (
            .AXLEN_W (AXLEN_W),
            .AW (AW),
            .DW (DW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP),
            .CMD_SIZE_W(CMD_SIZE_W),
            .CMD_UW (CMD_UW) 
) u_icb2axi_aw (
            .icb_cmd_valid (icb_cmd_valid_raw),
            .icb_cmd_ready (icb_cmd_ready_raw),
            .icb_cmd_addr (icb_cmd_addr), 
            .icb_cmd_xlen(icb_cmd_xlen),
            .icb_cmd_xburst(icb_cmd_xburst),
            .icb_cmd_modes (icb_cmd_modes ),
            .icb_cmd_dmode (icb_cmd_dmode ),
            .icb_cmd_attri (icb_cmd_attri ),
            .icb_cmd_read (icb_cmd_read), 
            .icb_cmd_wdata (icb_cmd_wdata),
            .icb_cmd_wmask (icb_cmd_wmask),
            .icb_cmd_beat (icb_cmd_beat),
            .icb_cmd_lock (icb_cmd_lock),
            .icb_cmd_excl (icb_cmd_excl),
            .icb_cmd_size (icb_cmd_size),
            .icb_cmd_usr (icb_cmd_usr),
            .axi_awready (axi_awready),
            .axi_awvalid (axi_awvalid),
            .axi_awaddr (axi_awaddr),
            .axi_awlen (axi_awlen),
            .axi_awsize (axi_awsize),
            .axi_awburst (axi_awburst),
            .axi_awlock (axi_awlock),
            .axi_awcache (axi_awcache),
            .axi_awprot (axi_awprot),
            .axi_awuser (axi_awuser),
            .axi_wready (axi_wready),
            .axi_wvalid (axi_wvalid),
            .axi_wdata (axi_wdata),
            .axi_wstrb (axi_wstrb),
            .axi_wlast (axi_wlast),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .clk (clk),
            .rst_n (rst_n)
  );
  e603_subsys_gnrl_ficb2axi_b # (
            .AW (AW),
            .DW (DW),
            .RSP_UW (RSP_UW),
        .PAYLOAD_NORST(PAYLOAD_NORST),
            .RATIO_FIFO_DP(RATIO_FIFO_DP) 
   ) u_icb2axi_b(
            .wrsp_burst_fifo_o_vld (wrsp_burst_fifo_o_vld),
            .icb_wrsp_valid (icb_rsp_valid),
            .icb_wrsp_ready (icb_rsp_ready),
            .icb_wrsp_err (icb_rsp_err),
            .icb_wrsp_excl_ok (icb_rsp_excl_ok),
            .icb_wrsp_usr (icb_rsp_usr),
            .axi_bready (axi_bready),
            .axi_bvalid (axi_bvalid),
            .axi_bresp (axi_bresp),
            .axi_buser (axi_buser),
            .axi_bus_clk_en (axi_bus_clk_en),
            .icb_clk_en (icb_clk_en),
            .wrsp_xlen  (wrsp_xlen),
            .wrsp_last  (wrsp_last),
            .clk (clk),
            .rst_n (rst_n)
  );
  assign icb2axi_write_pend_active = wrsp_burst_fifo_o_vld | axi_wvalid | axi_awvalid;
endmodule
module e603_subsys_gnrl_ficb2axi_read_async # (
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter OUTS_CNT_W = 4,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 1,
  parameter ASYNC_FIFO_DP = 6,
  parameter ASYNC_FIFO_DP_PTR_W = 3,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  output                        icb2axi_read_async_icb_active,
  output                        icb2axi_read_async_axi_active,
  output                        icb2axi_read_pend_active,
  input                         axi_arready,
  output                        axi_arvalid,
  output [AW-1:0]               axi_araddr,
  output [7:0]                  axi_arlen,
  output [CMD_SIZE_W-1:0]                  axi_arsize,
  output [1:0]                  axi_arburst,
  output                        axi_arlock,
  output [3:0]                  axi_arcache,
  output [2:0]                  axi_arprot,
  output [CMD_UW-1:0]            axi_aruser,
  output                        axi_rready,
  input                         axi_rvalid,
  input [DW-1:0]                axi_rdata,
  input [RSP_UW-1:0]             axi_ruser,
  input [1:0]                   axi_rresp,
  input                         axi_rlast,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [7:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]            icb_rsp_usr,
  input  async_axi_clk,
  input  async_axi_rst_n,
  input  icb_clk,
  input  icb_rst_n
  );
  wire i_icb_reset_flag_r;
e603_subsys_gnrl_dffrs #(1) reset_flag_dffrs (1'b0, i_icb_reset_flag_r, icb_clk, icb_rst_n);// VPP_NO_REG_PARSE
  wire i_icb_cmd_valid;
  wire i_icb_cmd_ready;
  assign i_icb_cmd_valid = (~i_icb_reset_flag_r) & icb_cmd_valid;
  assign icb_cmd_ready   = (~i_icb_reset_flag_r) & i_icb_cmd_ready;
  wire                        icb2axi_arready;
  wire                        icb2axi_arvalid;
  wire [AW-1:0]               icb2axi_araddr;
  wire [7:0]                  icb2axi_arlen;
  wire [CMD_SIZE_W-1:0]                  icb2axi_arsize;
  wire [1:0]                  icb2axi_arburst;
  wire                        icb2axi_arlock;
  wire [3:0]                  icb2axi_arcache;
  wire [2:0]                  icb2axi_arprot;
  wire [CMD_UW-1:0]           icb2axi_aruser;
  localparam AR_PACK_W = (AW+8+CMD_SIZE_W+2+1+4+3+CMD_UW) 
          ;
  wire [AR_PACK_W-1:0] ar_fifo_i_dat = {
                              icb2axi_araddr,
                              icb2axi_arlen,
                              icb2axi_arsize,
                              icb2axi_arburst,
                              icb2axi_arlock,
                              icb2axi_arcache,
                              icb2axi_arprot,
                              icb2axi_aruser 
                                 };
  wire [AR_PACK_W-1:0] ar_fifo_o_dat;
  assign {
                              axi_araddr,
                              axi_arlen,
                              axi_arsize,
                              axi_arburst,
                              axi_arlock,
                              axi_arcache,
                              axi_arprot,
                              axi_aruser
                                } = ar_fifo_o_dat;
  wire                        icb2axi_rready;
  wire                        icb2axi_rvalid;
  wire[DW-1:0]                icb2axi_rdata;
  wire[RSP_UW-1:0]            icb2axi_ruser;
  wire[1:0]                   icb2axi_rresp;
  wire                        icb2axi_rlast;
  localparam R_PACK_W = (1+2+DW+RSP_UW);
  wire [R_PACK_W-1:0] r_fifo_i_dat = {
                              axi_rdata,
                              axi_ruser,
                              axi_rresp,
                              axi_rlast 
                                 };
  wire [R_PACK_W-1:0] r_fifo_o_dat;
  assign {
                              icb2axi_rdata,
                              icb2axi_ruser,
                              icb2axi_rresp,
                              icb2axi_rlast 
                                 } = r_fifo_o_dat;
wire i_icb2axi_read_pend_active;
 e603_subsys_gnrl_ficb2axi_read # (
            .AW (AW),
            .DW (DW),
            .OUTS_CNT_W(OUTS_CNT_W),
            .RATIO_FIFO_DP(0),
            .CMD_UW (CMD_UW),
            .RSP_UW (RSP_UW)
   ) u_icb2axi_read(
            .icb2axi_read_pend_active(i_icb2axi_read_pend_active),
            .icb_cmd_valid    (i_icb_cmd_valid),
            .icb_cmd_ready    (i_icb_cmd_ready),
            .icb_cmd_addr     (icb_cmd_addr), 
            .icb_cmd_sel      (icb_cmd_sel), 
            .icb_cmd_xlen     (icb_cmd_xlen),
            .icb_cmd_xburst   (icb_cmd_xburst),
            .icb_cmd_modes    (icb_cmd_modes ),
            .icb_cmd_dmode    (icb_cmd_dmode ),
            .icb_cmd_attri    (icb_cmd_attri ),
            .icb_cmd_read     (icb_cmd_read), 
            .icb_cmd_wdata    (icb_cmd_wdata),
            .icb_cmd_wmask    (icb_cmd_wmask),
            .icb_cmd_beat     (icb_cmd_beat),
            .icb_cmd_lock     (icb_cmd_lock),
            .icb_cmd_excl     (icb_cmd_excl),
            .icb_cmd_size     (icb_cmd_size),
            .icb_cmd_usr      (icb_cmd_usr),
            .icb_rsp_valid   (icb_rsp_valid),
            .icb_rsp_ready   (icb_rsp_ready),
            .icb_rsp_rdata   (icb_rsp_rdata),
            .icb_rsp_usr     (icb_rsp_usr),
            .icb_rsp_err     (icb_rsp_err),
            .icb_rsp_excl_ok (icb_rsp_excl_ok),
            .axi_arready (icb2axi_arready),
            .axi_arvalid (icb2axi_arvalid),
            .axi_araddr  (icb2axi_araddr),
            .axi_arlen   (icb2axi_arlen),
            .axi_arsize  (icb2axi_arsize),
            .axi_arburst (icb2axi_arburst),
            .axi_arlock  (icb2axi_arlock),
            .axi_arcache (icb2axi_arcache),
            .axi_arprot  (icb2axi_arprot),
            .axi_aruser  (icb2axi_aruser),
            .axi_rready (icb2axi_rready),
            .axi_rvalid (icb2axi_rvalid),
            .axi_rdata  (icb2axi_rdata),
            .axi_ruser  (icb2axi_ruser),
            .axi_rresp  (icb2axi_rresp),
            .axi_rlast  (icb2axi_rlast),
            .axi_bus_clk_en (1'b1),
            .icb_clk_en (1'b1),
            .clk   (icb_clk),
            .rst_n (icb_rst_n) 
  );
  wire ar_async_i_active;
  wire ar_async_o_active;
  wire r_async_i_active;
  wire r_async_o_active;
  e603_subsys_gnrl_cdc_fifo # (
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (AR_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_ar(
    .i_clk   (icb_clk),
    .i_rst_n (icb_rst_n),
    .o_clk   (async_axi_clk),
    .o_rst_n (async_axi_rst_n),
    .i_vld    (icb2axi_arvalid),
    .i_rdy    (icb2axi_arready),
    .i_dat    (ar_fifo_i_dat),
    .i_cdc_fifo_active(ar_async_i_active),
    .o_cdc_fifo_active(ar_async_o_active),
    .o_vld    (axi_arvalid),
    .o_rdy    (axi_arready),
    .o_dat    (ar_fifo_o_dat )
  );
  e603_subsys_gnrl_cdc_fifo # (
    .DP(ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (R_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_r(
    .o_clk   (icb_clk),
    .o_rst_n (icb_rst_n), 
    .i_clk   (async_axi_clk),
    .i_rst_n (async_axi_rst_n),
    .i_vld   (axi_rvalid),
    .i_rdy   (axi_rready),
    .i_dat   (r_fifo_i_dat ),
    .i_cdc_fifo_active(r_async_i_active),
    .o_cdc_fifo_active(r_async_o_active),
    .o_vld  (icb2axi_rvalid),
    .o_rdy  (icb2axi_rready),
    .o_dat  (r_fifo_o_dat )
  );
  wire axi2axi_async_i_active = ar_async_i_active | r_async_o_active ;
  wire axi2axi_async_o_active = ar_async_o_active | r_async_i_active ;
  assign icb2axi_read_async_icb_active = i_icb2axi_read_pend_active | axi2axi_async_i_active;
  assign icb2axi_read_async_axi_active = axi2axi_async_o_active;
  assign icb2axi_read_pend_active = icb2axi_read_async_icb_active;
endmodule
module e603_subsys_gnrl_ficb2axi_write_async # (
  parameter OUTS_CNT_W =2,
  parameter OUTS_FIFO_DP =4,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 1,
  parameter ASYNC_FIFO_DP = 6,
  parameter ASYNC_FIFO_DP_PTR_W = 3,
  parameter CMD_UW = 1,
  parameter RSP_UW = 1
  ) (
  output                        icb2axi_write_async_icb_active,
  output                        icb2axi_write_async_axi_active,
  output                        icb2axi_write_pend_active,
  input                         axi_awready,
  output                        axi_awvalid,
  output [AW-1:0]               axi_awaddr,
  output [7:0]                  axi_awlen,
  output [CMD_SIZE_W-1:0]                  axi_awsize,
  output [1:0]                  axi_awburst,
  output                        axi_awlock,
  output [3:0]                  axi_awcache,
  output [2:0]                  axi_awprot,
  output [CMD_UW-1:0]            axi_awuser, 
  input                         axi_wready,
  output                        axi_wvalid,
  output [DW-1:0]               axi_wdata,
  output [DW/8-1:0]               axi_wstrb,
  output                        axi_wlast,
  output                         axi_bready,
  input                          axi_bvalid,
  input [RSP_UW-1:0]              axi_buser,
  input [1:0]                    axi_bresp,
  input                         icb_cmd_sel,
  input                         icb_cmd_valid,
  output                        icb_cmd_ready,
  input [AW-1:0]                icb_cmd_addr, 
  input                         icb_cmd_read, 
  input [DW-1:0]                icb_cmd_wdata,
  input [DW/8-1:0]                icb_cmd_wmask,
  input [CMD_UW-1:0]             icb_cmd_usr,
  input [1:0]                   icb_cmd_beat,
  input                         icb_cmd_lock,
  input                         icb_cmd_excl,
  input [CMD_SIZE_W-1:0]                   icb_cmd_size,
  input [7:0]                   icb_cmd_xlen,
  input [1:0]                   icb_cmd_xburst,
  input [1:0]                   icb_cmd_modes,
  input                         icb_cmd_dmode,
  input [2:0]                   icb_cmd_attri,
  output                        icb_rsp_valid,
  input                         icb_rsp_ready,
  output                        icb_rsp_err  ,
  output                        icb_rsp_excl_ok,
  output [DW-1:0]               icb_rsp_rdata,
  output [RSP_UW-1:0]            icb_rsp_usr,
  input  async_axi_clk,
  input  async_axi_rst_n,
  input  icb_clk,
  input  icb_rst_n
  );
  wire i_icb_reset_flag_r;
e603_subsys_gnrl_dffrs #(1) reset_flag_dffrs (1'b0, i_icb_reset_flag_r, icb_clk, icb_rst_n);// VPP_NO_REG_PARSE
  wire i_icb_cmd_valid;
  wire i_icb_cmd_ready;
  assign i_icb_cmd_valid = (~i_icb_reset_flag_r) & icb_cmd_valid;
  assign icb_cmd_ready   = (~i_icb_reset_flag_r) & i_icb_cmd_ready;
  wire aw_async_i_active;
  wire aw_async_o_active;
  wire w_async_i_active ;
  wire w_async_o_active ;
  wire b_async_o_active ;
  wire b_async_i_active ;
  wire axi2axi_async_i_active = aw_async_i_active | w_async_i_active | b_async_o_active ;
  wire axi2axi_async_o_active = aw_async_o_active | w_async_o_active | b_async_i_active ;
  wire                        icb2axi_awready;
  wire                        icb2axi_awvalid;
  wire [AW-1:0]               icb2axi_awaddr;
  wire [7:0]                  icb2axi_awlen;
  wire [CMD_SIZE_W-1:0]                  icb2axi_awsize;
  wire [1:0]                  icb2axi_awburst;
  wire                        icb2axi_awlock;
  wire [3:0]                  icb2axi_awcache;
  wire [2:0]                  icb2axi_awprot;
  wire [CMD_UW-1:0]           icb2axi_awuser;
  localparam AW_PACK_W = (AW+8+CMD_SIZE_W+2+1+4+3+CMD_UW) 
                       ;
  wire [AW_PACK_W-1:0] aw_fifo_i_dat = {
                              icb2axi_awaddr,
                              icb2axi_awlen,
                              icb2axi_awsize,
                              icb2axi_awburst,
                              icb2axi_awlock,
                              icb2axi_awcache,
                              icb2axi_awprot,
                              icb2axi_awuser 
                                 };
  wire [AW_PACK_W-1:0] aw_fifo_o_dat;
  assign {
                              axi_awaddr,
                              axi_awlen,
                              axi_awsize,
                              axi_awburst,
                              axi_awlock,
                              axi_awcache,
                              axi_awprot,
                              axi_awuser
                                } = aw_fifo_o_dat;
  e603_subsys_gnrl_cdc_fifo # (
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (AW_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_aw(
    .i_clk   (icb_clk),
    .i_rst_n (icb_rst_n),
    .o_clk   (async_axi_clk),
    .o_rst_n (async_axi_rst_n),
    .i_vld    (icb2axi_awvalid),
    .i_rdy    (icb2axi_awready),
    .i_dat    (aw_fifo_i_dat),
    .i_cdc_fifo_active(aw_async_i_active),
    .o_cdc_fifo_active(aw_async_o_active),
    .o_vld    (axi_awvalid),
    .o_rdy    (axi_awready),
    .o_dat    (aw_fifo_o_dat )
  );
  wire                        icb2axi_wready;
  wire                        icb2axi_wvalid;
  wire [DW-1:0]               icb2axi_wdata;
  wire [DW/8-1:0]             icb2axi_wstrb;
  wire                        icb2axi_wlast;
  localparam W_PACK_W = (DW+(DW/8)+1);
  wire [W_PACK_W-1:0] w_fifo_i_dat = {
                              icb2axi_wdata,
                              icb2axi_wstrb,
                              icb2axi_wlast 
                                 };
  wire [W_PACK_W-1:0] w_fifo_o_dat;
  assign {
                              axi_wdata,
                              axi_wstrb,
                              axi_wlast 
                                } = w_fifo_o_dat;
  e603_subsys_gnrl_cdc_fifo # (
    .DP     (ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (W_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_w(
    .i_clk   (icb_clk),
    .i_rst_n (icb_rst_n), 
    .o_clk   (async_axi_clk),
    .o_rst_n (async_axi_rst_n),
    .i_vld    (icb2axi_wvalid),
    .i_rdy    (icb2axi_wready),
    .i_dat    (w_fifo_i_dat),
    .i_cdc_fifo_active(w_async_i_active),
    .o_cdc_fifo_active(w_async_o_active),
    .o_vld    (axi_wvalid),
    .o_rdy    (axi_wready),
    .o_dat    (w_fifo_o_dat )
  );
  wire icb2axi_bvalid;
  wire icb2axi_bready;
  wire [RSP_UW-1:0] icb2axi_buser;
  wire [1:0]        icb2axi_bresp;
  localparam B_PACK_W = (2+RSP_UW);
  wire [B_PACK_W-1:0] b_fifo_i_dat = {
                                 axi_buser,
                                 axi_bresp 
                                 };
  wire [B_PACK_W-1:0] b_fifo_o_dat;
  assign {
                              icb2axi_buser,
                              icb2axi_bresp 
                                 } = b_fifo_o_dat;
  e603_subsys_gnrl_cdc_fifo # (
    .DP(ASYNC_FIFO_DP),
    .DP_PTR_W     (ASYNC_FIFO_DP_PTR_W),
    .DW     (B_PACK_W),
    .SYNC_DP(SYNC_DP)
  ) u_cdc_fifo_b(
    .o_clk   (icb_clk),
    .o_rst_n (icb_rst_n), 
    .i_clk   (async_axi_clk),
    .i_rst_n (async_axi_rst_n),
    .i_vld   (axi_bvalid),
    .i_rdy   (axi_bready),
    .i_dat   (b_fifo_i_dat ),
    .i_cdc_fifo_active(b_async_i_active),
    .o_cdc_fifo_active(b_async_o_active),
    .o_vld  (icb2axi_bvalid),
    .o_rdy  (icb2axi_bready),
    .o_dat  (b_fifo_o_dat )
  );
  wire i_icb2axi_write_pend_active;
 e603_subsys_gnrl_ficb2axi_write # (
            .AW (AW),
            .DW (DW),
            .RATIO_FIFO_DP(0),
            .OUTS_CNT_W  (OUTS_CNT_W ),
            .OUTS_FIFO_DP  (OUTS_FIFO_DP ),
            .CMD_UW (CMD_UW),
            .RSP_UW (RSP_UW)
   ) u_icb2axi_write(
            .icb2axi_write_pend_active(i_icb2axi_write_pend_active),
            .icb_cmd_valid   (i_icb_cmd_valid),
            .icb_cmd_ready   (i_icb_cmd_ready),
            .icb_cmd_addr    (icb_cmd_addr), 
            .icb_cmd_sel     (icb_cmd_sel), 
            .icb_cmd_xlen    (icb_cmd_xlen),
            .icb_cmd_xburst  (icb_cmd_xburst),
            .icb_cmd_modes   (icb_cmd_modes ),
            .icb_cmd_dmode   (icb_cmd_dmode ),
            .icb_cmd_attri   (icb_cmd_attri ),
            .icb_cmd_read    (icb_cmd_read), 
            .icb_cmd_wdata   (icb_cmd_wdata),
            .icb_cmd_wmask   (icb_cmd_wmask),
            .icb_cmd_beat    (icb_cmd_beat),
            .icb_cmd_lock    (icb_cmd_lock),
            .icb_cmd_excl    (icb_cmd_excl),
            .icb_cmd_size    (icb_cmd_size),
            .icb_cmd_usr     (icb_cmd_usr),
            .icb_rsp_valid   (icb_rsp_valid),
            .icb_rsp_ready   (icb_rsp_ready),
            .icb_rsp_rdata   (icb_rsp_rdata),
            .icb_rsp_usr     (icb_rsp_usr),
            .icb_rsp_err     (icb_rsp_err),
            .icb_rsp_excl_ok (icb_rsp_excl_ok),
            .axi_awready (icb2axi_awready ),
            .axi_awvalid (icb2axi_awvalid ),
            .axi_awaddr  (icb2axi_awaddr  ),
            .axi_awlen   (icb2axi_awlen   ),
            .axi_awsize  (icb2axi_awsize  ),
            .axi_awburst (icb2axi_awburst ),
            .axi_awlock  (icb2axi_awlock  ),
            .axi_awcache (icb2axi_awcache ),
            .axi_awprot  (icb2axi_awprot  ),
            .axi_awuser  (icb2axi_awuser  ),
            .axi_wready  (icb2axi_wready  ),
            .axi_wvalid  (icb2axi_wvalid  ),
            .axi_wdata   (icb2axi_wdata   ),
            .axi_wstrb   (icb2axi_wstrb   ),
            .axi_wlast   (icb2axi_wlast   ),
            .axi_bready  (icb2axi_bready  ),
            .axi_bvalid  (icb2axi_bvalid  ),
            .axi_buser   (icb2axi_buser   ),
            .axi_bresp   (icb2axi_bresp   ),
            .axi_bus_clk_en (1'b1),
            .icb_clk_en (1'b1),
            .clk   (icb_clk),
            .rst_n (icb_rst_n)
  );
  assign icb2axi_write_async_icb_active = i_icb2axi_write_pend_active | axi2axi_async_i_active;
  assign icb2axi_write_async_axi_active = axi2axi_async_o_active;
  assign icb2axi_write_pend_active = icb2axi_write_async_icb_active;
endmodule
`include "global.v"
module  e603_subsys_gnrl_axi2ficb_write # (
  parameter PAYLOAD_NORST = 0,
  parameter ALLOW_FIX_BURST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           axi_awready,
  input                            axi_awvalid,
  input [ID_W-1:0]        axi_awid,
  input [AW-1:0]      axi_awaddr,
  input [7:0]                      axi_awlen,
  input [CMD_SIZE_W-1:0]                      axi_awsize,
  input [1:0]                      axi_awburst,
  input                            axi_awlock,
  input [3:0]                      axi_awcache,
  input [2:0]                      axi_awprot,
  input [USR_W-1:0]          axi_awuser, 
  output                           axi_wready,
  input                            axi_wvalid,
  input [DW-1:0]           axi_wdata,
  input [MW-1:0]        axi_wstrb,
  input                            axi_wlast,
  input                            axi_bready,
  output                           axi_bvalid,
  output [USR_W-1:0]          axi_buser, 
  output [ID_W-1:0]       axi_bid,
  output [1:0]                     axi_bresp,
  output                           icb_wcmd_sel,
  output                           icb_wcmd_valid,
  input                            icb_wcmd_ready,
  output [AW-1:0]                  icb_wcmd_addr,
  output                           icb_wcmd_read, 
  output [DW-1:0]                  icb_wcmd_wdata,
  output [MW-1:0]                  icb_wcmd_wmask,
  output [1:0]                     icb_wcmd_beat,
  output                           icb_wcmd_lock,
  output                           icb_wcmd_excl,
  output [CMD_SIZE_W-1:0]         icb_wcmd_size,
  output [7:0]                     icb_wcmd_xlen,
  output [1:0]                     icb_wcmd_xburst,
  output [1:0]                     icb_wcmd_modes,
  output                           icb_wcmd_dmode,
  output [2:0]                     icb_wcmd_attri,
  output [USR_W-1:0]               icb_wcmd_usr,
  input                            icb_wrsp_valid,
  output                           icb_wrsp_ready,
  input                            icb_wrsp_err,
  input                            icb_wrsp_excl_ok,
  input  [USR_W-1:0]               icb_wrsp_usr,
  input                            axi_bus_clk_en,
  input                            icb_clk_en,
  output                           axi2icb_write_active,
  input  clk,
  input  rst_n
  );
  wire axi_awready_raw;
  wire axi_awvalid_raw;
  wire axi_wready_raw;
  wire axi_wvalid_raw;
  assign axi_awvalid_raw = (~reset_flag_r) & axi_awvalid    ;
  assign axi_awready     = (~reset_flag_r) & axi_awready_raw;
  assign axi_wvalid_raw  = (~reset_flag_r) & axi_wvalid    ;
  assign axi_wready      = (~reset_flag_r) & axi_wready_raw;
  assign icb_wcmd_lock = 1'b0;
    localparam AXI_AW_BUF_PACK = ID_W+AW+8+CMD_SIZE_W+2+1+3+4+USR_W;
    wire [AXI_AW_BUF_PACK-1:0] i_axi_aw_pack = {
                                             axi_awid    ,  
                                             axi_awaddr  ,
                                             axi_awlen   ,
                                             axi_awsize  ,
                                             axi_awburst ,
                                             axi_awlock  ,
                                             axi_awcache ,
                                             axi_awprot  ,
                                             axi_awuser   
                                            };
    wire [ID_W-1:0]    axi_buf_o_awid    ; 
    wire [AW-1:0]  axi_buf_o_awaddr  ; 
    wire [7:0]                  axi_buf_o_awlen   ; 
    wire [CMD_SIZE_W-1:0]                  axi_buf_o_awsize  ; 
    wire [1:0]                  axi_buf_o_awburst ; 
    wire                        axi_buf_o_awlock  ; 
    wire [3:0]                  axi_buf_o_awcache ; 
    wire [2:0]                  axi_buf_o_awprot  ; 
    wire [USR_W-1:0]      axi_buf_o_awuser  ; 
    wire [AXI_AW_BUF_PACK-1:0] o_axi_aw_pack ;
    assign  { 
              axi_buf_o_awid    , 
              axi_buf_o_awaddr  , 
              axi_buf_o_awlen   , 
              axi_buf_o_awsize  , 
              axi_buf_o_awburst , 
              axi_buf_o_awlock  , 
              axi_buf_o_awcache , 
              axi_buf_o_awprot  , 
              axi_buf_o_awuser    
            } = o_axi_aw_pack ;
    wire axi_buf_o_awvalid ;    
    wire axi_buf_o_awready ; 
    wire axi_o_awbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_AW_BUF_PACK)
    ) u_axi_aw_fifo(
    .i_clk_en(axi_bus_clk_en), 
    .i_vld(axi_awvalid_raw  ), 
    .i_rdy(axi_awready_raw  ), 
    .i_dat(i_axi_aw_pack),
    .o_clk_en(icb_clk_en),
    .o_vld(axi_buf_o_awvalid), 
    .o_rdy(axi_buf_o_awready), 
    .o_dat(o_axi_aw_pack    ),
    .o_fifo_active(axi_o_awbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
    localparam AXI_W_BUF_PACK = DW+MW+1;
    wire [AXI_W_BUF_PACK-1:0] i_axi_w_pack = {
                                             axi_wdata      , 
                                             axi_wstrb      , 
                                             axi_wlast        
                                            };
    wire [DW-1:0]       axi_buf_o_wdata  ; 
    wire [MW-1:0]    axi_buf_o_wstrb  ; 
    wire                        axi_buf_o_wlast  ; 
    wire [AXI_W_BUF_PACK-1:0] o_axi_w_pack ;
    assign  { 
              axi_buf_o_wdata  , 
              axi_buf_o_wstrb  , 
              axi_buf_o_wlast    
            } = o_axi_w_pack ;
    wire axi_buf_o_wvalid ;    
    wire axi_buf_o_wready ; 
    wire axi_o_wbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_W_BUF_PACK)
    ) u_axi_w_fifo(
    .i_clk_en(axi_bus_clk_en),
    .i_vld(axi_wvalid_raw  ), 
    .i_rdy(axi_wready_raw  ), 
    .i_dat(i_axi_w_pack),
    .o_clk_en(icb_clk_en),
    .o_vld(axi_buf_o_wvalid), 
    .o_rdy(axi_buf_o_wready), 
    .o_dat(o_axi_w_pack    ),
    .o_fifo_active(axi_o_wbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire axi_buf_o_awready_pos;
  wire axi_buf_o_awvalid_pos;
  wire write_id_fifo_rdy;
  assign axi_buf_o_awready     = write_id_fifo_rdy & axi_buf_o_awready_pos;
  assign axi_buf_o_awvalid_pos = write_id_fifo_rdy & axi_buf_o_awvalid    ;
  e603_subsys_gnrl_axi2ficb_aw # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W),
    .USR_W (USR_W)
  ) u_aw_axi2icb(
    .axi_awready  (axi_buf_o_awready_pos ),
    .axi_awvalid  (axi_buf_o_awvalid_pos & icb_clk_en ),
    .axi_awid     (axi_buf_o_awid    ),
    .axi_awaddr   (axi_buf_o_awaddr  ),
    .axi_awlen    (axi_buf_o_awlen   ),
    .axi_awsize   (axi_buf_o_awsize  ),
    .axi_awburst  (axi_buf_o_awburst ),
    .axi_awlock   (axi_buf_o_awlock  ),
    .axi_awcache  (axi_buf_o_awcache ),
    .axi_awprot   (axi_buf_o_awprot  ),
    .axi_awuser   (axi_buf_o_awuser),
    .axi_wready   (axi_buf_o_wready),
    .axi_wvalid   (axi_buf_o_wvalid & icb_clk_en),
    .axi_wdata    (axi_buf_o_wdata ),
    .axi_wstrb    (axi_buf_o_wstrb ),
    .axi_wlast    (axi_buf_o_wlast ),
    .icb_wcmd_sel (icb_wcmd_sel),
    .icb_wcmd_valid (icb_wcmd_valid),
    .icb_wcmd_ready (icb_wcmd_ready & icb_clk_en),
    .icb_wcmd_addr  (icb_wcmd_addr ), 
    .icb_wcmd_read  (icb_wcmd_read ), 
    .icb_wcmd_wdata (icb_wcmd_wdata),
    .icb_wcmd_wmask (icb_wcmd_wmask),
    .icb_wcmd_beat  (icb_wcmd_beat ),
    .icb_wcmd_lock  (              ), 
    .icb_wcmd_excl  (icb_wcmd_excl ),
    .icb_wcmd_size  (icb_wcmd_size ),
    .icb_wcmd_xlen    (icb_wcmd_xlen   ),
    .icb_wcmd_xburst  (icb_wcmd_xburst ),
    .icb_wcmd_modes   (icb_wcmd_modes  ),
    .icb_wcmd_dmode   (icb_wcmd_dmode  ),
    .icb_wcmd_attri   (icb_wcmd_attri  ),
    .icb_wcmd_usr   (icb_wcmd_usr  ), 
    .clk (clk),
    .rst_n (rst_n)
  );
    localparam AXI_B_BUF_PACK = ID_W+2+USR_W;
    wire [USR_W-1:0]   axi_buf_i_buser    ; 
    wire [ID_W-1:0]    axi_buf_i_bid    ; 
    wire [1:0]                  axi_buf_i_bresp  ; 
    wire [AXI_B_BUF_PACK-1:0] i_axi_b_pack = {
                                             axi_buf_i_buser  ,  
                                             axi_buf_i_bid  ,  
                                             axi_buf_i_bresp        
                                            };
    wire [AXI_B_BUF_PACK-1:0] o_axi_b_pack ;
    assign  { 
              axi_buser    , 
              axi_bid    , 
              axi_bresp    
            } = o_axi_b_pack ;
    wire axi_buf_i_bvalid ;    
    wire axi_buf_i_bready ; 
    wire axi_o_bbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_B_BUF_PACK)
    ) u_axi_b_fifo(
    .i_clk_en(icb_clk_en),
    .i_vld(axi_buf_i_bvalid), 
    .i_rdy(axi_buf_i_bready), 
    .i_dat(i_axi_b_pack    ),
    .o_clk_en(axi_bus_clk_en),
    .o_vld(axi_bvalid  ), 
    .o_rdy(axi_bready  ), 
    .o_dat(o_axi_b_pack),
    .o_fifo_active(axi_o_bbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire write_id_fifo_active;
  wire [7:0] wrsp_xlen;
  wire  wrsp_burst;
  e603_subsys_gnrl_axi2ficb_b # (
    .USR_W (USR_W),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W)
  ) u_b_axi2icb(
    .icb_wrsp_ready   (icb_wrsp_ready  ),
    .icb_wrsp_valid   (icb_wrsp_valid  & icb_clk_en),
    .icb_wrsp_err     (icb_wrsp_err    ),
    .icb_wrsp_usr     (icb_wrsp_usr    ),
    .icb_wrsp_excl_ok (icb_wrsp_excl_ok),
    .axi_bready       (axi_buf_i_bready & icb_clk_en),
    .axi_bvalid       (axi_buf_i_bvalid),
    .axi_bresp        (axi_buf_i_bresp ),
    .axi_buser        (axi_buf_i_buser ),
    .axi_bid          (axi_buf_i_bid   ), 
    .wrsp_xlen_vld  (write_id_fifo_active),
    .wrsp_xlen  (wrsp_xlen),
    .wrsp_burst (wrsp_burst),
    .clk (clk),
    .rst_n (rst_n)
  );
  wire wcmd_burst = (~(axi_buf_o_awlen == 8'b0)) ;
  wire [7:0] wcmd_xlen  = axi_buf_o_awlen;
  localparam WRSP_FIFO_PACK = 1+8+ID_W;
  e603_subsys_gnrl_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .CUT_READY (1),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
        .DW  (WRSP_FIFO_PACK)
  ) u_wrsp_fifo (
        .i_vld(axi_buf_o_awvalid && axi_buf_o_awready & icb_clk_en),
        .i_rdy(write_id_fifo_rdy),
        .i_dat({wcmd_burst,wcmd_xlen, axi_buf_o_awid}),
        .o_vld(write_id_fifo_active),
        .o_rdy(axi_buf_i_bvalid && axi_buf_i_bready & icb_clk_en ),  
        .o_dat({wrsp_burst,wrsp_xlen, 
                      axi_buf_i_bid
                      }),  
        .clk  (clk),
        .rst_n(rst_n)
  );
   assign axi2icb_write_active = axi_o_awbusy | axi_o_wbusy | axi_o_bbusy 
                               | write_id_fifo_active
                               ;
endmodule
module  e603_subsys_gnrl_axi2ficb_read # (
  parameter PAYLOAD_NORST = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           axi_arready,
  input                            axi_arvalid,
  input [ID_W-1:0]        axi_arid,
  input [AW-1:0]      axi_araddr,
  input [7:0]                      axi_arlen,
  input [CMD_SIZE_W-1:0]                      axi_arsize,
  input [1:0]                      axi_arburst,
  input                            axi_arlock,
  input [3:0]                      axi_arcache,
  input [2:0]                      axi_arprot,
  input [USR_W-1:0]          axi_aruser,
  input                            axi_rready,
  output                           axi_rvalid,
  output [ID_W-1:0]       axi_rid,
  output [DW-1:0]          axi_rdata,
  output [1:0]                     axi_rresp,
  output                           axi_rlast,
  output [USR_W-1:0]          axi_ruser,
  output                           icb_rcmd_sel ,
  output                           icb_rcmd_valid ,
  input                            icb_rcmd_ready ,
  output [AW-1:0]                  icb_rcmd_addr  ,
  output                           icb_rcmd_read  ,
  output [DW-1:0]                  icb_rcmd_wdata ,
  output [MW-1:0]                  icb_rcmd_wmask ,
  output [1:0]                     icb_rcmd_beat  ,
  output                           icb_rcmd_excl  ,             
  output [CMD_SIZE_W-1:0]         icb_rcmd_size  ,
  output [7:0]                     icb_rcmd_xlen,
  output [1:0]                     icb_rcmd_xburst,
  output [1:0]                     icb_rcmd_modes,
  output                           icb_rcmd_dmode,
  output [2:0]                     icb_rcmd_attri,
  output [USR_W-1:0]               icb_rcmd_usr   ,
  output                           icb_rrsp_ready  , 
  input                            icb_rrsp_valid  , 
  input [DW-1:0]                   icb_rrsp_rdata  , 
  input                            icb_rrsp_err    , 
  input                            icb_rrsp_excl_ok, 
  input [USR_W-1:0]                icb_rrsp_usr   ,
  input                            axi_bus_clk_en,
  input                            icb_clk_en,
  output                           axi2icb_read_active,
  input clk  ,
  input rst_n  
  );
  wire axi_arvalid_raw;
  wire axi_arready_raw;
  assign axi_arvalid_raw = (~reset_flag_r) & axi_arvalid;
  assign axi_arready     = (~reset_flag_r) & axi_arready_raw;
    localparam AXI_AR_BUF_PACK = ID_W+AW+8+CMD_SIZE_W+2+1+3+4+USR_W;
    wire [AXI_AR_BUF_PACK-1:0] i_axi_ar_pack = {
                                             axi_arid    ,  
                                             axi_araddr  ,
                                             axi_arlen   ,
                                             axi_arsize  ,
                                             axi_arburst ,
                                             axi_arlock  ,
                                             axi_arcache ,
                                             axi_arprot  ,
                                             axi_aruser   
                                            };
    wire [ID_W-1:0]    axi_buf_o_arid    ; 
    wire [AW-1:0]  axi_buf_o_araddr  ; 
    wire [7:0]                  axi_buf_o_arlen   ; 
    wire [CMD_SIZE_W-1:0]                  axi_buf_o_arsize  ; 
    wire [1:0]                  axi_buf_o_arburst ; 
    wire                        axi_buf_o_arlock  ; 
    wire [3:0]                  axi_buf_o_arcache ; 
    wire [2:0]                  axi_buf_o_arprot  ; 
    wire [USR_W-1:0]      axi_buf_o_aruser  ; 
    wire [AXI_AR_BUF_PACK-1:0] o_axi_ar_pack ;
    assign  { 
              axi_buf_o_arid    , 
              axi_buf_o_araddr  , 
              axi_buf_o_arlen   , 
              axi_buf_o_arsize  , 
              axi_buf_o_arburst , 
              axi_buf_o_arlock  , 
              axi_buf_o_arcache , 
              axi_buf_o_arprot  , 
              axi_buf_o_aruser    
            } = o_axi_ar_pack ;
    wire axi_buf_o_arvalid ;    
    wire axi_buf_o_arready ; 
    wire axi_o_arbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_AR_BUF_PACK)
    ) u_axi_ar_fifo(
    .i_clk_en(axi_bus_clk_en), 
    .i_vld(axi_arvalid_raw      ), 
    .i_rdy(axi_arready_raw      ), 
    .i_dat(i_axi_ar_pack    ),
    .o_clk_en(icb_clk_en), 
    .o_vld(axi_buf_o_arvalid), 
    .o_rdy(axi_buf_o_arready), 
    .o_dat(o_axi_ar_pack    ),
    .o_fifo_active(axi_o_arbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire axi_buf_o_arready_pos;
  wire axi_buf_o_arvalid_pos;
  wire read_id_fifo_rdy;
  assign axi_buf_o_arready     = read_id_fifo_rdy & axi_buf_o_arready_pos;
  assign axi_buf_o_arvalid_pos = read_id_fifo_rdy & axi_buf_o_arvalid;
  e603_subsys_gnrl_axi2ficb_ar # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W),
    .USR_W (USR_W)  
  ) u_ar_axi2icb(
     .axi_arready  (axi_buf_o_arready_pos ),
     .axi_arvalid  (axi_buf_o_arvalid_pos & icb_clk_en ),
     .axi_arid     (axi_buf_o_arid    ),
     .axi_araddr   (axi_buf_o_araddr  ),
     .axi_arlen    (axi_buf_o_arlen   ),
     .axi_arsize   (axi_buf_o_arsize  ),
     .axi_arburst  (axi_buf_o_arburst ),
     .axi_arlock   (axi_buf_o_arlock  ),
     .axi_arcache  (axi_buf_o_arcache ),
     .axi_arprot   (axi_buf_o_arprot  ),
     .axi_aruser   (axi_buf_o_aruser), 
     .icb_rcmd_sel   (icb_rcmd_sel),
     .icb_rcmd_valid (icb_rcmd_valid),
     .icb_rcmd_ready (icb_rcmd_ready & icb_clk_en),
     .icb_rcmd_addr  (icb_rcmd_addr ), 
     .icb_rcmd_read  (icb_rcmd_read ), 
     .icb_rcmd_wdata (icb_rcmd_wdata),
     .icb_rcmd_wmask (icb_rcmd_wmask),
     .icb_rcmd_beat  (icb_rcmd_beat ),
     .icb_rcmd_lock  (              ), 
     .icb_rcmd_excl  (icb_rcmd_excl ),
     .icb_rcmd_size  (icb_rcmd_size ),
     .icb_rcmd_xlen    (icb_rcmd_xlen   ),
     .icb_rcmd_xburst  (icb_rcmd_xburst ),
     .icb_rcmd_modes   (icb_rcmd_modes  ),
     .icb_rcmd_dmode   (icb_rcmd_dmode  ),
     .icb_rcmd_attri   (icb_rcmd_attri  ),
     .icb_rcmd_usr   (icb_rcmd_usr  ),
     .clk   (clk),
     .rst_n (rst_n)
  );
    localparam AXI_R_BUF_PACK = USR_W+ID_W+DW+2+1;
    wire [USR_W-1:0]    axi_buf_i_ruser    ; 
    wire [ID_W-1:0]    axi_buf_i_rid    ; 
    wire [ID_W-1:0]    axi_rid_from_fifo    ; 
    wire [DW-1:0]       axi_buf_i_rdata  ; 
    wire [1:0]                  axi_buf_i_rresp  ; 
    wire                        axi_buf_i_rlast  ; 
    wire [AXI_R_BUF_PACK-1:0] i_axi_r_pack = {
                                             axi_buf_i_ruser    ,
                                             axi_buf_i_rid    ,
                                             axi_buf_i_rdata  ,
                                             axi_buf_i_rresp  ,
                                             axi_buf_i_rlast   
                                            };
    wire [AXI_R_BUF_PACK-1:0] o_axi_r_pack ;
    assign  { 
              axi_ruser        ,  
              axi_rid        ,  
              axi_rdata      ,  
              axi_rresp      ,  
              axi_rlast         
            } = o_axi_r_pack ;
    wire axi_buf_i_rvalid ;    
    wire axi_buf_i_rready ; 
    wire axi_o_rbusy ; 
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_R_BUF_PACK)
    ) u_axi_r_fifo(
    .i_clk_en(icb_clk_en),
    .i_vld(axi_buf_i_rvalid), 
    .i_rdy(axi_buf_i_rready), 
    .i_dat(i_axi_r_pack    ),
    .o_clk_en(axi_bus_clk_en),
    .o_vld(axi_rvalid  ), 
    .o_rdy(axi_rready  ), 
    .o_dat(o_axi_r_pack),
    .o_fifo_active(axi_o_rbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
  wire [7:0] rrsp_xlen ;
  wire  rrsp_burst;
  wire read_id_fifo_active;
  e603_subsys_gnrl_axi2ficb_r # (
    .USR_W (USR_W),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ID_W (ID_W)
  ) u_axi2icb_r(
    .icb_rrsp_ready   (icb_rrsp_ready  ),
    .icb_rrsp_valid   (icb_rrsp_valid  & icb_clk_en  ),
    .icb_rrsp_rdata   (icb_rrsp_rdata  ),
    .icb_rrsp_usr     (icb_rrsp_usr    ),
    .icb_rrsp_err     (icb_rrsp_err    ),
    .icb_rrsp_excl_ok (icb_rrsp_excl_ok),
    .axi_rready       (axi_buf_i_rready & icb_clk_en),
    .axi_rvalid       (axi_buf_i_rvalid),
    .axi_rid          (axi_buf_i_rid   ),
    .axi_rid_from_fifo(axi_rid_from_fifo),
    .axi_ruser        (axi_buf_i_ruser ),
    .axi_rdata        (axi_buf_i_rdata ),
    .axi_rresp        (axi_buf_i_rresp ),
    .axi_rlast        (axi_buf_i_rlast ),
    .rrsp_xlen_vld    (read_id_fifo_active),
    .rrsp_xlen        (rrsp_xlen     ),
    .rrsp_burst       (rrsp_burst    ),
    .clk   (clk          ),
    .rst_n (rst_n)
  );
  wire rcmd_burst = (~(axi_buf_o_arlen == 8'b0)) ;
  wire [7:0] rcmd_xlen  = axi_buf_o_arlen;
  localparam RRSP_FIFO_PACK = 1+8+ID_W;
  e603_subsys_gnrl_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
        .CUT_READY (1),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM), 
        .DW  (RRSP_FIFO_PACK)
  ) u_rrsp_fifo (
        .i_vld(axi_buf_o_arvalid && axi_buf_o_arready  & icb_clk_en), 
        .i_rdy(read_id_fifo_rdy),
        .o_vld(read_id_fifo_active),
        .o_rdy(axi_buf_i_rvalid && axi_buf_i_rready && axi_buf_i_rlast  & icb_clk_en ),  
        .i_dat({rcmd_burst,rcmd_xlen, axi_buf_o_arid}),
        .o_dat({rrsp_burst,rrsp_xlen, axi_rid_from_fifo }),  
        .clk  (clk),
        .rst_n(rst_n)
  );
  assign axi2icb_read_active = axi_o_arbusy | axi_o_rbusy 
                             | read_id_fifo_active
                             ;
endmodule
module  e603_subsys_gnrl_axi2ficb_ar # (
  parameter PAYLOAD_NORST = 0,
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ID_W = 4, 
  parameter USR_W = 1
) (
  output                         axi_arready,
  input                          axi_arvalid,
  input [ID_W-1:0]               axi_arid,
  input [AW-1:0]                 axi_araddr,
  input [7:0]                    axi_arlen,
  input [CMD_SIZE_W-1:0]                    axi_arsize,
  input [1:0]                    axi_arburst,
  input                          axi_arlock,
  input [3:0]                    axi_arcache,
  input [2:0]                    axi_arprot,
  input [USR_W-1:0]              axi_aruser,
  output                         icb_rcmd_valid,
  input                          icb_rcmd_ready,
  output [AW-1:0]                icb_rcmd_addr, 
  output                         icb_rcmd_read, 
  output [DW-1:0]                icb_rcmd_wdata,
  output [MW-1:0]                icb_rcmd_wmask,
  output [1:0]                   icb_rcmd_beat,
  output                         icb_rcmd_lock,
  output                         icb_rcmd_excl,
  output [CMD_SIZE_W-1:0]       icb_rcmd_size,
  output [USR_W-1:0]             icb_rcmd_usr,
  output                         icb_rcmd_sel,
  output [7:0]                   icb_rcmd_xlen,
  output [1:0]                   icb_rcmd_xburst,
  output [1:0]                   icb_rcmd_modes,
  output                         icb_rcmd_dmode,
  output [2:0]                   icb_rcmd_attri,
  input                         clk,
  input                         rst_n
  );
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_nxt;
  wire       burst_cnt_ena;
  wire       rcmd_burst;
  wire       rcmd_burst_r;
  wire axi_arlock_buf;
  wire [CMD_SIZE_W-1:0] axi_arsize_buf;
  wire [1:0] axi_arburst_buf;
  wire [7:0] axi_arlen_buf;
  wire [2:0] axi_arprot_buf ;
  wire [3:0] axi_arcache_buf;
  wire [USR_W-1:0] axi_aruser_buf;
  wire [ID_W-1:0] axi_arid_buf;
  wire [AW-1:0] axi_araddr_buf;
  wire buf_wr_en;
  assign rcmd_burst = axi_arvalid  & (~(axi_arlen == 8'b0)) ;
  wire burst_first = (burst_cnt_r == 8'b0);
  assign rcmd_burst_r = ~burst_first;
  assign burst_cnt_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_last = (burst_cnt_r == axi_arlen_buf) & (~burst_first);
  assign burst_cnt_ena = (rcmd_burst || rcmd_burst_r) && icb_rcmd_valid && icb_rcmd_ready;
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign buf_wr_en = rcmd_burst && icb_rcmd_valid && icb_rcmd_ready && burst_first;
  generate
  if(PAYLOAD_NORST == 1) begin: payload_norst 
e603_subsys_gnrl_dffl  #(1) arlock_dffl  ( buf_wr_en, axi_arlock, axi_arlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(CMD_SIZE_W) arsize_dffl  ( buf_wr_en, axi_arsize, axi_arsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(8) arlen_dffl  ( buf_wr_en, axi_arlen, axi_arlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2) arburst_dffl  ( buf_wr_en, axi_arburst, axi_arburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(USR_W) aruser_dffl  ( buf_wr_en, axi_aruser, axi_aruser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(3) arprot_dffl   ( buf_wr_en, axi_arprot,  axi_arprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(4) arcache_dffl  ( buf_wr_en, axi_arcache, axi_arcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(ID_W) arid_dffl  ( buf_wr_en, axi_arid, axi_arid_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: payload_rst
e603_subsys_gnrl_dfflr #(1) arlock_dfflr ( buf_wr_en, axi_arlock, axi_arlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(CMD_SIZE_W) arsize_dfflr ( buf_wr_en, axi_arsize, axi_arsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(8) arlen_dfflr ( buf_wr_en, axi_arlen, axi_arlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(2) arburst_dfflr ( buf_wr_en, axi_arburst, axi_arburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(USR_W) aruser_dfflr ( buf_wr_en, axi_aruser, axi_aruser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(3) arprot_dfflr  ( buf_wr_en, axi_arprot,  axi_arprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(4) arcache_dfflr ( buf_wr_en, axi_arcache, axi_arcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(ID_W) arid_dfflr ( buf_wr_en, axi_arid, axi_arid_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  assign axi_arready   = icb_rcmd_ready && (!rcmd_burst_r);
  assign icb_rcmd_valid   = axi_arvalid  || rcmd_burst_r;
  wire icb_rcmd_read_tmp    = 1'b1; 
  assign icb_rcmd_read = icb_rcmd_read_tmp;
  assign icb_rcmd_wdata   = {DW{1'b0}};
  assign icb_rcmd_wmask   = {MW{1'b0}};
  wire icb_rcmd_lock_tmp    = 1'b0; 
  assign icb_rcmd_lock    = icb_rcmd_lock_tmp;
  wire icb_rcmd_excl_tmp    = rcmd_burst_r ? axi_arlock_buf : axi_arlock;
  assign icb_rcmd_excl = icb_rcmd_excl_tmp;
  wire [CMD_SIZE_W-1:0] icb_rcmd_size_tmp;
  assign icb_rcmd_size_tmp    = rcmd_burst_r ? axi_arsize_buf[CMD_SIZE_W-1:0] : axi_arsize[CMD_SIZE_W-1:0];
  assign icb_rcmd_size = icb_rcmd_size_tmp;
  wire icb_rcmd_fxed;
  wire icb_rcmd_incr;
  wire icb_rcmd_wrap;
  wire axi_araddr_ena = burst_cnt_ena;
  wire [AW-1:0] icb_rcmd_addr_mask = ({AW{1'b1}} << icb_rcmd_size);
  wire [AW-1:0] icb_rcmd_addr_algned = (icb_rcmd_addr_mask & icb_rcmd_addr);
  wire [12-1:0] axi_araddr_incr_size = (icb_rcmd_addr_algned[11:0] + (12'b1 << icb_rcmd_size));
  wire [12-1:0] axi_araddr_wrap_mask = ((~{8'b0,icb_rcmd_xlen[3:0]}) << icb_rcmd_size);
  wire [12-1:0] axi_araddr_incr_wrap = (axi_araddr_incr_size & (~axi_araddr_wrap_mask)) | (icb_rcmd_addr[11:0] & axi_araddr_wrap_mask);
  wire [AW-1:0] axi_araddr_nxt = icb_rcmd_fxed ? icb_rcmd_addr : 
                                 icb_rcmd_wrap ? {icb_rcmd_addr[AW-1:12],axi_araddr_incr_wrap} :
                                                 {icb_rcmd_addr[AW-1:12],axi_araddr_incr_size};
  generate
  if(PAYLOAD_NORST == 1) begin: araddr_payload_norst 
e603_subsys_gnrl_dffl  #(AW) araddr_dffl  ( axi_araddr_ena, axi_araddr_nxt, axi_araddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: araddr_payload_rst
e603_subsys_gnrl_dfflr #(AW) araddr_dfflr ( axi_araddr_ena, axi_araddr_nxt, axi_araddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  wire icb_rcmd_xlen_eq3  = (icb_rcmd_xlen == 8'd3) ;
  wire icb_rcmd_xlen_eq7  = (icb_rcmd_xlen == 8'd7) ;
  wire icb_rcmd_xlen_eq15 = (icb_rcmd_xlen == 8'd15);
  assign icb_rcmd_fxed = (icb_rcmd_xburst == 2'b00);
  assign icb_rcmd_incr = (icb_rcmd_xburst == 2'b01);
  assign icb_rcmd_wrap = (icb_rcmd_xburst == 2'b10);
  wire icb_rcmd_xburst_fixed;
  wire [1:0] icb_rcmd_beat_tmp;
  assign icb_rcmd_beat_tmp  = icb_rcmd_xburst_fixed          ? 2'b00 :
                          ( rcmd_burst && !rcmd_burst_r) ? 2'b01 : 
                          (burst_last)                   ? 2'b10 :
                                                           2'b00 ;
  assign icb_rcmd_beat = icb_rcmd_beat_tmp;
  wire [AW-1:0] icb_rcmd_addr_raw; 
  assign icb_rcmd_addr_raw  = (!rcmd_burst_r) ? axi_araddr :
                          axi_araddr_buf ; 
  assign icb_rcmd_usr   = rcmd_burst_r ? axi_aruser_buf : axi_aruser;
  wire [2:0] icb_rcmd_arprot  = rcmd_burst_r ? axi_arprot_buf  : axi_arprot;
  wire [3:0] icb_rcmd_arcache = rcmd_burst_r ? axi_arcache_buf : axi_arcache;
  wire [7:0] icb_rcmd_arlen   = rcmd_burst_r ? axi_arlen_buf   : axi_arlen;
  wire [AW-1:0] icb_rcmd_addr_tmp;
  assign icb_rcmd_addr_tmp  = icb_rcmd_addr_raw;
  assign icb_rcmd_addr = icb_rcmd_addr_tmp; 
  wire icb_rcmd_nonalloc = (icb_rcmd_arcache == 4'b1011);
  wire icb_rcmd_device = icb_rcmd_nonalloc | (icb_rcmd_arcache == 4'b0000) | (icb_rcmd_arcache == 4'b0001);
  wire icb_rcmd_cacheb = (icb_rcmd_arcache == 4'b1111) | (icb_rcmd_arcache == 4'b0111) | (icb_rcmd_arcache == 4'b1011);
  wire icb_rcmd_nc     = icb_rcmd_nonalloc | ((~icb_rcmd_device) & (~icb_rcmd_cacheb));
  wire icb_rcmd_mmode = icb_rcmd_arprot[0];
  wire icb_rcmd_hmode = 1'b0;
  wire icb_rcmd_smode = 1'b0;
  wire icb_rcmd_ifu   = icb_rcmd_arprot[2];
  assign icb_rcmd_sel  = icb_rcmd_valid;
  wire [1:0] icb_rcmd_modes_tmp;
  assign icb_rcmd_modes_tmp = icb_rcmd_mmode ? 2'd0 : icb_rcmd_hmode ? 2'd1 : icb_rcmd_smode ? 2'd2 : 2'd3;
  assign icb_rcmd_modes = icb_rcmd_modes_tmp;
  wire icb_rcmd_dmode_tmp = 1'b0;
  assign icb_rcmd_dmode = icb_rcmd_dmode_tmp;
  wire [2:0] icb_rcmd_attri_tmp;
  assign icb_rcmd_attri_tmp[0] = icb_rcmd_ifu   ;
  assign icb_rcmd_attri_tmp[1] = icb_rcmd_device;
  assign icb_rcmd_attri_tmp[2] = icb_rcmd_nc    ;
  assign icb_rcmd_attri = icb_rcmd_attri_tmp;
  wire [7:0] icb_rcmd_xlen_tmp;
  assign icb_rcmd_xlen_tmp = icb_rcmd_xburst_fixed ? 8'd0 : icb_rcmd_arlen;
  assign icb_rcmd_xlen = icb_rcmd_xlen_tmp;
  generate 
      if(ALLOW_FIX_BURST == 1) begin: allow_fix_burst_gen
  assign icb_rcmd_xburst_fixed = 1'b0;
      end
      else begin: disallow_fix_burst_gen
  assign icb_rcmd_xburst_fixed = (icb_rcmd_xburst == 2'b00);
      end
  endgenerate
  wire [1:0] icb_rcmd_xburst_tmp; 
  assign icb_rcmd_xburst_tmp = rcmd_burst_r ? axi_arburst_buf : axi_arburst;
  assign icb_rcmd_xburst = icb_rcmd_xburst_tmp;
endmodule
module  e603_subsys_gnrl_axi2ficb_aw # (
  parameter PAYLOAD_NORST = 0,
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  output                         axi_awready,
  input                          axi_awvalid,
  input [ID_W-1:0]               axi_awid,
  input [AW-1:0]                 axi_awaddr,
  input [7:0]                    axi_awlen,
  input [CMD_SIZE_W-1:0]                    axi_awsize,
  input [1:0]                    axi_awburst,
  input                          axi_awlock,
  input [3:0]                    axi_awcache,
  input [2:0]                    axi_awprot,
  input [USR_W-1:0]              axi_awuser,
  output                         axi_wready,
  input                          axi_wvalid,
  input [DW-1:0]                 axi_wdata,
  input [MW-1:0]                 axi_wstrb,
  input                          axi_wlast,
  output                         icb_wcmd_valid,
  input                          icb_wcmd_ready,
  output [AW-1:0]                icb_wcmd_addr, 
  output                         icb_wcmd_read, 
  output [DW-1:0]                icb_wcmd_wdata,
  output [MW-1:0]                icb_wcmd_wmask,
  output [1:0]                   icb_wcmd_beat,
  output                         icb_wcmd_lock,
  output                         icb_wcmd_excl,
  output [CMD_SIZE_W-1:0]       icb_wcmd_size,
  output [USR_W-1:0]             icb_wcmd_usr,
  output                         icb_wcmd_sel,
  output [7:0]                   icb_wcmd_xlen,
  output [1:0]                   icb_wcmd_xburst,
  output [1:0]                   icb_wcmd_modes,
  output                         icb_wcmd_dmode,
  output [2:0]                   icb_wcmd_attri,
  input                         clk,
  input                         rst_n
  );
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_nxt;
  wire       burst_cnt_ena;
  wire       wcmd_burst;
  wire       wcmd_burst_r;
  wire axi_awlock_buf;
  wire [CMD_SIZE_W-1:0] axi_awsize_buf;
  wire [1:0] axi_awburst_buf;
  wire [7:0] axi_awlen_buf;
  wire [USR_W-1:0] axi_awuser_buf;
  wire [AW-1:0] axi_awaddr_buf;
  wire [2:0] axi_awprot_buf ;
  wire [3:0] axi_awcache_buf;
  wire buf_wr_en;
  assign wcmd_burst = axi_awvalid  & (~(axi_awlen == 8'b0)) ;
  wire burst_first = (burst_cnt_r == 8'b0);
  assign wcmd_burst_r = ~burst_first;
  assign burst_cnt_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_last = (burst_cnt_r == axi_awlen_buf)& (~burst_first);
  assign burst_cnt_ena = (wcmd_burst || wcmd_burst_r) && icb_wcmd_valid && icb_wcmd_ready;
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign buf_wr_en = wcmd_burst && icb_wcmd_valid && icb_wcmd_ready && burst_first;
  generate
  if(PAYLOAD_NORST == 1) begin: payload_norst 
e603_subsys_gnrl_dffl  #(1) awlock_dffl  ( buf_wr_en, axi_awlock, axi_awlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(CMD_SIZE_W) awsize_dffl  ( buf_wr_en, axi_awsize, axi_awsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(8) awlen_dffl  ( buf_wr_en, axi_awlen, axi_awlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(2) awburst_dffl  ( buf_wr_en, axi_awburst, axi_awburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(USR_W) awuser_dffl  ( buf_wr_en, axi_awuser, axi_awuser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(3) awprot_dffl   ( buf_wr_en, axi_awprot,  axi_awprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dffl  #(4) awcache_dffl  ( buf_wr_en, axi_awcache, axi_awcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: payload_rst
e603_subsys_gnrl_dfflr #(1) awlock_dfflr ( buf_wr_en, axi_awlock, axi_awlock_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(CMD_SIZE_W) awsize_dfflr ( buf_wr_en, axi_awsize, axi_awsize_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(8) awlen_dfflr ( buf_wr_en, axi_awlen, axi_awlen_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(2) awburst_dfflr ( buf_wr_en, axi_awburst, axi_awburst_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(USR_W) awuser_dfflr ( buf_wr_en, axi_awuser, axi_awuser_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(3) awprot_dfflr  ( buf_wr_en, axi_awprot,  axi_awprot_buf, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(4) awcache_dfflr ( buf_wr_en, axi_awcache, axi_awcache_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  wire icb_wcmd_read_tmp; 
  assign icb_wcmd_read_tmp    = 1'b0; 
  assign icb_wcmd_read = icb_wcmd_read_tmp;
  wire [DW-1:0] icb_wcmd_wdata_tmp;
  wire [MW-1:0] icb_wcmd_wmask_tmp;
  assign icb_wcmd_wdata_tmp   = axi_wdata;
  assign icb_wcmd_wmask_tmp   = axi_wstrb;
  assign icb_wcmd_wdata = icb_wcmd_wdata_tmp;
  assign icb_wcmd_wmask = icb_wcmd_wmask_tmp;
  wire [CMD_SIZE_W-1:0] icb_wcmd_size_tmp;
  wire icb_wcmd_lock_tmp    = 1'b0;
  assign icb_wcmd_lock = icb_wcmd_lock_tmp;
  wire icb_wcmd_excl_tmp    = wcmd_burst_r ? axi_awlock_buf : axi_awlock;
  assign icb_wcmd_excl = icb_wcmd_excl_tmp;
  assign icb_wcmd_size_tmp    = wcmd_burst_r ? axi_awsize_buf[CMD_SIZE_W-1:0] : axi_awsize[CMD_SIZE_W-1:0];
  assign icb_wcmd_size    = icb_wcmd_size_tmp;
  assign axi_awready   = icb_wcmd_ready && (!wcmd_burst_r) && axi_wvalid;
  assign axi_wready    = icb_wcmd_ready && (wcmd_burst_r || axi_awvalid);
  assign icb_wcmd_valid   = (axi_awvalid || wcmd_burst_r) && axi_wvalid ;
  wire icb_wcmd_fxed;
  wire icb_wcmd_incr;
  wire icb_wcmd_wrap;
  wire axi_awaddr_ena = burst_cnt_ena;
  wire [AW-1:0] icb_wcmd_addr_mask = ({AW{1'b1}} << icb_wcmd_size);
  wire [AW-1:0] icb_wcmd_addr_algned = (icb_wcmd_addr_mask & icb_wcmd_addr);
  wire [12-1:0] axi_awaddr_incr_size = (icb_wcmd_addr_algned[11:0] + (12'b1 << icb_wcmd_size));
  wire [12-1:0] axi_awaddr_wrap_mask = ((~{8'b0,icb_wcmd_xlen[3:0]}) << icb_wcmd_size);
  wire [12-1:0] axi_awaddr_incr_wrap = (axi_awaddr_incr_size & (~axi_awaddr_wrap_mask)) | (icb_wcmd_addr[11:0] & axi_awaddr_wrap_mask);
  wire [AW-1:0] axi_awaddr_nxt = icb_wcmd_fxed ? icb_wcmd_addr : 
                                 icb_wcmd_wrap ? {icb_wcmd_addr[AW-1:12],axi_awaddr_incr_wrap} :
                                                 {icb_wcmd_addr[AW-1:12],axi_awaddr_incr_size};
    generate
  if(PAYLOAD_NORST == 1) begin: awaddr_payload_norst 
e603_subsys_gnrl_dffl  #(AW) awaddr_dffl  ( axi_awaddr_ena, axi_awaddr_nxt, axi_awaddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  else begin: awaddr_payload_rst
e603_subsys_gnrl_dfflr #(AW) awaddr_dfflr ( axi_awaddr_ena, axi_awaddr_nxt, axi_awaddr_buf, clk, rst_n);// VPP_NO_REG_PARSE
  end
  endgenerate
  wire icb_wcmd_xlen_eq3  = (icb_wcmd_xlen == 8'd3) ;
  wire icb_wcmd_xlen_eq7  = (icb_wcmd_xlen == 8'd7) ;
  wire icb_wcmd_xlen_eq15 = (icb_wcmd_xlen == 8'd15);
  assign icb_wcmd_fxed = (icb_wcmd_xburst == 2'b00);
  assign icb_wcmd_incr = (icb_wcmd_xburst == 2'b01);
  assign icb_wcmd_wrap = (icb_wcmd_xburst == 2'b10);
  wire icb_wcmd_xburst_fixed;
  wire [1:0] icb_wcmd_beat_tmp;
  assign icb_wcmd_beat_tmp  = icb_wcmd_xburst_fixed          ? 
                                        2'b00 :
                          ( wcmd_burst && !wcmd_burst_r) ? 2'b01 : 
                          (burst_last)                   ? 2'b10 :
                                                           2'b00 ;
  assign icb_wcmd_beat  = icb_wcmd_beat_tmp;
  wire [AW-1:0] icb_wcmd_addr_raw; 
  assign icb_wcmd_addr_raw  = (!wcmd_burst_r) ? axi_awaddr :
                          axi_awaddr_buf ; 
  assign icb_wcmd_usr   = wcmd_burst_r ? axi_awuser_buf : axi_awuser;
  wire [2:0] icb_wcmd_awprot  = wcmd_burst_r ? axi_awprot_buf  : axi_awprot;
  wire [3:0] icb_wcmd_awcache = wcmd_burst_r ? axi_awcache_buf : axi_awcache;
  wire [7:0] icb_wcmd_awlen   = wcmd_burst_r ? axi_awlen_buf   : axi_awlen;
  wire [AW-1:0] icb_wcmd_addr_tmp;
  assign icb_wcmd_addr_tmp  = icb_wcmd_addr_raw;
  assign icb_wcmd_addr = icb_wcmd_addr_tmp;  
  wire icb_wcmd_nonalloc = (icb_wcmd_awcache == 4'b0111);
  wire icb_wcmd_device = icb_wcmd_nonalloc | (icb_wcmd_awcache == 4'b0000) | (icb_wcmd_awcache == 4'b0001);
  wire icb_wcmd_cacheb = (icb_wcmd_awcache == 4'b1111) | (icb_wcmd_awcache == 4'b0111) | (icb_wcmd_awcache == 4'b1011);
  wire icb_wcmd_nc     = icb_wcmd_nonalloc | ((~icb_wcmd_device) & (~icb_wcmd_cacheb));
  wire icb_wcmd_mmode = icb_wcmd_awprot[0];
  wire icb_wcmd_hmode = 1'b0;
  wire icb_wcmd_smode = 1'b0;
  wire icb_wcmd_ifu   = icb_wcmd_awprot[2];
  assign icb_wcmd_sel  = icb_wcmd_valid;
  wire [1:0] icb_wcmd_modes_tmp = icb_wcmd_mmode ? 2'd0 : icb_wcmd_hmode ? 2'd1 : icb_wcmd_smode ? 2'd2 : 2'd3;
  assign icb_wcmd_modes = icb_wcmd_modes_tmp;
  wire icb_wcmd_dmode_tmp = 1'b0;
  wire [2:0] icb_wcmd_attri_tmp;
  assign icb_wcmd_dmode = icb_wcmd_dmode_tmp;
  assign icb_wcmd_attri_tmp[0] = icb_wcmd_ifu   ;
  assign icb_wcmd_attri_tmp[1] = icb_wcmd_device;
  assign icb_wcmd_attri_tmp[2] = icb_wcmd_nc    ;
  assign icb_wcmd_attri = icb_wcmd_attri_tmp;
  wire [1:0] icb_wcmd_xburst_tmp;
  assign icb_wcmd_xburst_tmp = wcmd_burst_r ? axi_awburst_buf : axi_awburst;
  assign icb_wcmd_xburst = icb_wcmd_xburst_tmp;
  wire [7:0] icb_wcmd_xlen_tmp;
  assign icb_wcmd_xlen_tmp = icb_wcmd_xburst_fixed ? 8'd0 : icb_wcmd_awlen;
  assign icb_wcmd_xlen = icb_wcmd_xlen_tmp;
  generate 
      if(ALLOW_FIX_BURST == 1) begin: allow_fix_burst_gen
  assign icb_wcmd_xburst_fixed = 1'b0;
      end
      else begin: disallow_fix_burst_gen
  assign icb_wcmd_xburst_fixed = (icb_wcmd_xburst == 2'b00);
      end
  endgenerate
endmodule
module  e603_subsys_gnrl_axi2ficb_r # (
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter USR_W = 4,
  parameter ID_W = 4
) (
  output                        icb_rrsp_ready,
  input                         icb_rrsp_valid,
  input [USR_W-1:0]             icb_rrsp_usr,
  input [DW-1:0]                icb_rrsp_rdata,
  input                         icb_rrsp_err,
  input                         icb_rrsp_excl_ok,
  input                         axi_rready,
  output                        axi_rvalid,
  output [USR_W-1:0]            axi_ruser,
  input  [ID_W-1:0]             axi_rid_from_fifo,
  output [ID_W-1:0]             axi_rid,
  output [DW-1:0]               axi_rdata,
  output [1:0]                  axi_rresp,
  output                        axi_rlast,
  input  [7:0]                  rrsp_xlen,
  input                         rrsp_burst,
  input                         rrsp_xlen_vld,
  input                         clk,
  input                         rst_n
  );
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_r_nxt;
  wire       burst_cnt_ena;
  wire burst_first = (burst_cnt_r == 8'd0);
  assign burst_cnt_r_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_last = (burst_cnt_r == rrsp_xlen) & (~burst_first);
  assign burst_cnt_ena = rrsp_burst && icb_rrsp_valid && icb_rrsp_ready;
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_r_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign icb_rrsp_ready   = rrsp_xlen_vld & axi_rready ;
  assign axi_rvalid       = rrsp_xlen_vld & icb_rrsp_valid ;
  wire [ID_W-1:0] axi_rid_tmp;
  assign axi_rid_tmp      = axi_rid_from_fifo;
  assign axi_rlast        = (!rrsp_burst) || (rrsp_burst && burst_last);
  wire [DW-1:0] axi_rdata_tmp;
  assign axi_rdata_tmp    = icb_rrsp_rdata;
  assign axi_ruser        = icb_rrsp_usr;
  assign axi_rresp        = {icb_rrsp_err,icb_rrsp_excl_ok};
  assign axi_rdata = axi_rdata_tmp;
  assign axi_rid = axi_rid_tmp; 
endmodule
module  e603_subsys_gnrl_axi2ficb_b # (
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter USR_W = 4,
  parameter ID_W = 4
) (
  output                        icb_wrsp_ready,
  input                         icb_wrsp_valid,
  input                         icb_wrsp_err,
  input                         icb_wrsp_excl_ok,
  input [USR_W-1:0]             icb_wrsp_usr,
  input                         axi_bready,
  output                        axi_bvalid,
  output [1:0]                  axi_bresp,
  input [ID_W-1:0]             axi_bid,
  output [USR_W-1:0]             axi_buser,
  input [7:0]                   wrsp_xlen,
  input                         wrsp_burst,
  input                         wrsp_xlen_vld,
  input                         clk,
  input                         rst_n
  );
  wire       burst_last;
  wire [7:0] burst_cnt_r;
  wire [7:0] burst_cnt_r_nxt;
  wire       burst_cnt_ena;
  assign burst_cnt_r_nxt = burst_last ? 8'b0 : (burst_cnt_r + 8'b1);
  assign burst_last = (burst_cnt_r == wrsp_xlen);
  assign burst_cnt_ena = wrsp_burst && icb_wrsp_valid && icb_wrsp_ready;
  assign icb_wrsp_ready   = ((wrsp_burst && !burst_last) || (axi_bready)) & wrsp_xlen_vld;
e603_subsys_gnrl_dfflr #(8) burst_cnt_dfflr (burst_cnt_ena, burst_cnt_r_nxt, burst_cnt_r, clk, rst_n);// VPP_NO_REG_PARSE
  assign axi_bvalid = (icb_wrsp_valid && (!wrsp_burst || (wrsp_burst && burst_last))) & wrsp_xlen_vld;
  wire [1:0]  axi_bresp_nxt;
  wire [1:0]  axi_bresp_buf;
  wire        axi_bresp_en;
  assign axi_bresp_en = wrsp_burst && icb_wrsp_valid && icb_wrsp_ready && !burst_last;
  assign axi_bresp_nxt = (burst_cnt_r == 0) ? {icb_wrsp_err,icb_wrsp_excl_ok}
                                             : (axi_bresp_buf | {icb_wrsp_err,icb_wrsp_excl_ok})
                                             ;
e603_subsys_gnrl_dfflr #(2) bresp_dfflr (axi_bresp_en, axi_bresp_nxt, axi_bresp_buf, clk, rst_n);// VPP_NO_REG_PARSE
  assign axi_bresp = ({2{wrsp_burst}} & axi_bresp_buf) | {icb_wrsp_err,icb_wrsp_excl_ok};
  assign axi_buser = icb_wrsp_usr;
endmodule
module  e603_subsys_gnrl_axi2ficb_read_async # (
  parameter ALLOW_FIX_BURST = 0,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 0,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input                            reset_flag_r,
  output                           axi_arready,
  input                            axi_arvalid,
  input [ID_W-1:0]                 axi_arid,
  input [AW-1:0]                   axi_araddr,
  input [7:0]                      axi_arlen,
  input [CMD_SIZE_W-1:0]                      axi_arsize,
  input [1:0]                      axi_arburst,
  input                            axi_arlock,
  input [3:0]                      axi_arcache,
  input [2:0]                      axi_arprot,
  input [USR_W-1:0]                axi_aruser,
  input                            axi_rready,
  output                           axi_rvalid,
  output [ID_W-1:0]                axi_rid,
  output [USR_W-1:0]               axi_ruser,
  output [DW-1:0]                  axi_rdata,
  output [1:0]                     axi_rresp,
  output                           axi_rlast,
  output                           icb_rcmd_sel   ,
  output                           icb_rcmd_valid ,
  input                            icb_rcmd_ready ,
  output [AW-1:0]                  icb_rcmd_addr  ,
  output                           icb_rcmd_read  ,
  output [DW-1:0]                  icb_rcmd_wdata ,
  output [MW-1:0]                  icb_rcmd_wmask ,
  output [1:0]                     icb_rcmd_beat  ,
  output                           icb_rcmd_excl  ,             
  output [CMD_SIZE_W-1:0]         icb_rcmd_size  ,
  output [7:0]                     icb_rcmd_xlen,
  output [1:0]                     icb_rcmd_xburst,
  output [1:0]                     icb_rcmd_modes,
  output                           icb_rcmd_dmode,
  output [2:0]                     icb_rcmd_attri,
  output [USR_W-1:0]               icb_rcmd_usr   ,
  output                           icb_rrsp_ready  , 
  input                            icb_rrsp_valid  , 
  input [DW-1:0]                   icb_rrsp_rdata  , 
  input [USR_W-1:0]                icb_rrsp_usr  , 
  input                            icb_rrsp_err    , 
  input                            icb_rrsp_excl_ok, 
  output                           axi2icb_read_axi_active,
  output                           axi2icb_read_icb_active,
  input icb_clk  ,
  input icb_rst_n,  
  input async_axi_clk  ,
  input async_axi_rst_n  
  );
  wire                           o_axi_arready;
  wire                           o_axi_arvalid;
  wire[ID_W-1:0]                 o_axi_arid;
  wire[AW-1:0]                   o_axi_araddr;
  wire[7:0]                      o_axi_arlen;
  wire[CMD_SIZE_W-1:0]                      o_axi_arsize;
  wire[1:0]                      o_axi_arburst;
  wire                           o_axi_arlock;
  wire[3:0]                      o_axi_arcache;
  wire[2:0]                      o_axi_arprot;
  wire[USR_W-1:0]                o_axi_aruser;
  wire                           o_axi_rready;
  wire                           o_axi_rvalid;
  wire [ID_W-1:0]                o_axi_rid;
  wire [USR_W-1:0]                o_axi_ruser;
  wire [DW-1:0]                  o_axi_rdata;
  wire [1:0]                     o_axi_rresp;
  wire                           o_axi_rlast;
  wire axi_buf_pipe_i_active;
  wire axi_buf_pipe_o_active;
  e603_subsys_gnrl_axi_buf_read # (
     .ASYNC (1),
     .SYNC_DP (SYNC_DP),
     .ASYNC_FIFO (ASYNC_FIFO),
     .ASYNC_FIFO_DP (ASYNC_FIFO_DP),
     .ASYNC_FIFO_DP_PTR_W (ASYNC_FIFO_DP_PTR_W),
     .RATIO_FIFO_DP(0),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW   (AW   ),
    .DW   (DW   ),
    .MW   (MW   ),
    .ID_W (ID_W ),
    .USR_W(USR_W) 
  ) u_axi_async_read(
    .reset_flag_r(reset_flag_r),
    .i_axi_arready        (axi_arready),
    .i_axi_arvalid        (axi_arvalid),
    .i_axi_arid           (axi_arid   ),
    .i_axi_araddr         (axi_araddr ),
    .i_axi_arlen          (axi_arlen  ),
    .i_axi_arsize         (axi_arsize ),
    .i_axi_arburst        (axi_arburst),
    .i_axi_arlock         (axi_arlock ),
    .i_axi_arcache        (axi_arcache),
    .i_axi_arprot         (axi_arprot ),
    .i_axi_aruser         (axi_aruser ),
    .i_axi_rready         (axi_rready ),
    .i_axi_rvalid         (axi_rvalid ),
    .i_axi_rid            (axi_rid    ),
    .i_axi_ruser          (axi_ruser    ),
    .i_axi_rdata          (axi_rdata  ),
    .i_axi_rresp          (axi_rresp  ),
    .i_axi_rlast          (axi_rlast  ),
    .o_axi_arready        (o_axi_arready),
    .o_axi_arvalid        (o_axi_arvalid),
    .o_axi_arid           (o_axi_arid   ),
    .o_axi_araddr         (o_axi_araddr ),
    .o_axi_arlen          (o_axi_arlen  ),
    .o_axi_arsize         (o_axi_arsize ),
    .o_axi_arburst        (o_axi_arburst),
    .o_axi_arlock         (o_axi_arlock ),
    .o_axi_arcache        (o_axi_arcache),
    .o_axi_arprot         (o_axi_arprot ),
    .o_axi_aruser         (o_axi_aruser ),
    .o_axi_rready         (o_axi_rready ),
    .o_axi_rvalid         (o_axi_rvalid ),
    .o_axi_rid            (o_axi_rid    ),
    .o_axi_ruser          (o_axi_ruser),
    .o_axi_rdata          (o_axi_rdata  ),
    .o_axi_rresp          (o_axi_rresp  ),
    .o_axi_rlast          (o_axi_rlast  ),
    .axi_buf_pipe_i_active  (axi_buf_pipe_i_active),
    .axi_buf_pipe_o_active  (axi_buf_pipe_o_active),
    .i_clk                (async_axi_clk  ),
    .i_rst_n              (async_axi_rst_n),
    .o_clk                (icb_clk  ),
    .o_rst_n              (icb_rst_n),
    .axi_bus_clk_en       (1'b1),
    .icb_clk_en           (1'b1),
    .clk                  (1'b0),
    .rst_n                (1'b0)  
  );
  wire o_axi2icb_read_active;
  e603_subsys_gnrl_axi2ficb_read # (
     .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
     .AW(AW),
     .DW(DW),
     .MW(MW),
     .RATIO_FIFO_DP(0),
     .FIFO_OUTS_NUM(FIFO_OUTS_NUM),
     .ID_W (ID_W),
     .USR_W (USR_W)
  ) u_axi2icb_read (
    .reset_flag_r    (1'b0),
    .axi_arready     (o_axi_arready ),
    .axi_arvalid     (o_axi_arvalid ),
    .axi_arid        (o_axi_arid    ),
    .axi_araddr      (o_axi_araddr  ),
    .axi_arlen       (o_axi_arlen   ),
    .axi_arsize      (o_axi_arsize  ),
    .axi_arburst     (o_axi_arburst ),
    .axi_arlock      (o_axi_arlock  ),
    .axi_arcache     (o_axi_arcache ),
    .axi_arprot      (o_axi_arprot  ),
    .axi_aruser      (o_axi_aruser  ),
    .axi_rready      (o_axi_rready   ),
    .axi_rvalid      (o_axi_rvalid   ),
    .axi_ruser       (o_axi_ruser    ),
    .axi_rid         (o_axi_rid      ),
    .axi_rdata       (o_axi_rdata    ),
    .axi_rresp       (o_axi_rresp    ),
    .axi_rlast       (o_axi_rlast    ),
    .icb_rcmd_sel    (icb_rcmd_sel    ),
    .icb_rcmd_valid  (icb_rcmd_valid  ),
    .icb_rcmd_ready  (icb_rcmd_ready  ),
    .icb_rcmd_addr   (icb_rcmd_addr   ),
    .icb_rcmd_read   (icb_rcmd_read   ),
    .icb_rcmd_wdata  (icb_rcmd_wdata  ),
    .icb_rcmd_wmask  (icb_rcmd_wmask  ),
    .icb_rcmd_beat   (icb_rcmd_beat   ),
    .icb_rcmd_excl   (icb_rcmd_excl   ),             
    .icb_rcmd_size   (icb_rcmd_size   ),
    .icb_rcmd_xlen   (icb_rcmd_xlen   ),
    .icb_rcmd_xburst (icb_rcmd_xburst ),
    .icb_rcmd_modes  (icb_rcmd_modes  ),
    .icb_rcmd_dmode  (icb_rcmd_dmode  ),
    .icb_rcmd_attri  (icb_rcmd_attri  ),
    .icb_rcmd_usr    (icb_rcmd_usr    ),
    .icb_rrsp_ready  (icb_rrsp_ready  ), 
    .icb_rrsp_valid  (icb_rrsp_valid  ), 
    .icb_rrsp_rdata  (icb_rrsp_rdata  ), 
    .icb_rrsp_err    (icb_rrsp_err    ), 
    .icb_rrsp_excl_ok(icb_rrsp_excl_ok), 
    .icb_rrsp_usr     (icb_rrsp_usr), 
    .axi_bus_clk_en  (1'b1),
    .icb_clk_en      (1'b1),
    .axi2icb_read_active  (o_axi2icb_read_active),
    .clk  (icb_clk  ),
    .rst_n(icb_rst_n)  
  );
  assign axi2icb_read_axi_active = axi_buf_pipe_i_active;
  assign axi2icb_read_icb_active = axi_buf_pipe_o_active | o_axi2icb_read_active;
endmodule
module  e603_subsys_gnrl_axi_buf_read # (
  parameter PAYLOAD_NORST = 0,
  parameter ASYNC = 0,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 0,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           i_axi_arready,
  input                            i_axi_arvalid,
  input [ID_W-1:0]                 i_axi_arid,
  input [AW-1:0]                   i_axi_araddr,
  input [AXLEN_W-1:0]                      i_axi_arlen,
  input [CMD_SIZE_W-1:0]                      i_axi_arsize,
  input [1:0]                      i_axi_arburst,
  input                            i_axi_arlock,
  input [3:0]                      i_axi_arcache,
  input [2:0]                      i_axi_arprot,
  input [USR_W-1:0]                i_axi_aruser,
  input                            i_axi_rready,
  output                           i_axi_rvalid,
  output [ID_W-1:0]                i_axi_rid,
  output [USR_W-1:0]               i_axi_ruser,
  output [DW-1:0]                  i_axi_rdata,
  output [1:0]                     i_axi_rresp,
  output                           i_axi_rlast,
  input                            o_axi_arready,
  output                           o_axi_arvalid,
  output[ID_W-1:0]                 o_axi_arid,
  output[AW-1:0]                   o_axi_araddr,
  output[AXLEN_W-1:0]                      o_axi_arlen,
  output[CMD_SIZE_W-1:0]                      o_axi_arsize,
  output[1:0]                      o_axi_arburst,
  output                           o_axi_arlock,
  output[3:0]                      o_axi_arcache,
  output[2:0]                      o_axi_arprot,
  output[USR_W-1:0]                o_axi_aruser,
  output                           o_axi_rready,
  input                            o_axi_rvalid,
  input  [ID_W-1:0]                o_axi_rid,
  input  [USR_W-1:0]               o_axi_ruser,
  input  [DW-1:0]                  o_axi_rdata,
  input  [1:0]                     o_axi_rresp,
  input                            o_axi_rlast,
  input                            axi_bus_clk_en,
  input                            icb_clk_en,
  output                           axi_buf_pipe_i_active,
  output                           axi_buf_pipe_o_active,
  input  i_clk,
  input  i_rst_n,
  input  o_clk,
  input  o_rst_n,
  input clk  ,
  input rst_n  
  );
  wire i_axi_arvalid_raw;
  wire i_axi_arready_raw;
  assign i_axi_arvalid_raw = (~reset_flag_r) & i_axi_arvalid;
  assign i_axi_arready     = (~reset_flag_r) & i_axi_arready_raw;
    localparam AXI_AR_BUF_PACK = ID_W+AW+AXLEN_W+CMD_SIZE_W+2+1+3+4+USR_W;
    wire [AXI_AR_BUF_PACK-1:0] i_axi_ar_pack = {
                                             i_axi_arid    ,  
                                             i_axi_araddr  ,
                                             i_axi_arlen   ,
                                             i_axi_arsize  ,
                                             i_axi_arburst ,
                                             i_axi_arlock  ,
                                             i_axi_arcache ,
                                             i_axi_arprot  ,
                                             i_axi_aruser   
                                            };
    wire [AXI_AR_BUF_PACK-1:0] o_axi_ar_pack ;
    assign  { 
              o_axi_arid    , 
              o_axi_araddr  , 
              o_axi_arlen   , 
              o_axi_arsize  , 
              o_axi_arburst , 
              o_axi_arlock  , 
              o_axi_arcache , 
              o_axi_arprot  , 
              o_axi_aruser    
            } = o_axi_ar_pack ;
    wire axi_i_arbusy ; 
    wire axi_o_arbusy ; 
    generate 
      if(ASYNC == 1) begin: ar_async_gen
        if(ASYNC_FIFO == 0) begin: ar_async_buf_gen
      e603_subsys_gnrl_cdc_buf
      # (
        .DW  (AXI_AR_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_ar_cdc_buf (
        .i_clk  (i_clk  ),
        .i_rst_n(i_rst_n),
        .i_vld(i_axi_arvalid_raw      ), 
        .i_rdy(i_axi_arready_raw      ), 
        .i_dat(i_axi_ar_pack    ),
        .i_cdc_buf_active(axi_i_arbusy), 
        .o_cdc_buf_active(axi_o_arbusy),
        .o_clk  (o_clk  ),
        .o_rst_n(o_rst_n),
        .o_vld(o_axi_arvalid), 
        .o_rdy(o_axi_arready), 
        .o_dat(o_axi_ar_pack    ) 
      );
       end
       else begin: ar_async_fifo_gen
      e603_subsys_gnrl_cdc_fifo
      # (
        .DP(ASYNC_FIFO_DP),
        .DP_PTR_W (ASYNC_FIFO_DP_PTR_W),
        .DW  (AXI_AR_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_ar_cdc_fifo (
        .i_clk  (i_clk  ),
        .i_rst_n(i_rst_n),
        .i_vld(i_axi_arvalid_raw      ), 
        .i_rdy(i_axi_arready_raw      ), 
        .i_dat(i_axi_ar_pack    ),
        .i_cdc_fifo_active(axi_i_arbusy), 
        .o_cdc_fifo_active(axi_o_arbusy),
        .o_clk  (o_clk  ),
        .o_rst_n(o_rst_n),
        .o_vld(o_axi_arvalid), 
        .o_rdy(o_axi_arready), 
        .o_dat(o_axi_ar_pack    ) 
      );
       end
      end
      else begin: ar_sync_gen
      assign axi_i_arbusy = i_axi_arvalid_raw;
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_AR_BUF_PACK)
    ) u_axi_ar_fifo(
    .i_clk_en(axi_bus_clk_en), 
    .i_vld(i_axi_arvalid_raw      ), 
    .i_rdy(i_axi_arready_raw      ), 
    .i_dat(i_axi_ar_pack    ),
    .o_clk_en(icb_clk_en), 
    .o_vld(o_axi_arvalid), 
    .o_rdy(o_axi_arready), 
    .o_dat(o_axi_ar_pack    ),
    .o_fifo_active(axi_o_arbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
      end
    endgenerate
    localparam AXI_R_BUF_PACK = USR_W + ID_W+DW+2+1;
    wire [AXI_R_BUF_PACK-1:0] i_axi_r_pack = {
                                             o_axi_ruser    ,
                                             o_axi_rid    ,
                                             o_axi_rdata  ,
                                             o_axi_rresp  ,
                                             o_axi_rlast   
                                            };
    wire [AXI_R_BUF_PACK-1:0] o_axi_r_pack ;
    assign  { 
              i_axi_ruser        ,  
              i_axi_rid        ,  
              i_axi_rdata      ,  
              i_axi_rresp      ,  
              i_axi_rlast         
            } = o_axi_r_pack ;
    wire axi_buf_i_rvalid ;    
    wire axi_buf_i_rready ; 
    wire axi_i_rbusy ; 
    wire axi_o_rbusy ; 
    generate 
      if(ASYNC == 1) begin: r_async_gen
        if(ASYNC_FIFO == 0) begin: r_async_buf_gen
      e603_subsys_gnrl_cdc_buf
      # (
        .DW  (AXI_R_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_r_cdc_buf (
        .i_clk  (o_clk  ),
        .i_rst_n(o_rst_n),
        .i_vld(o_axi_rvalid), 
        .i_rdy(o_axi_rready), 
        .i_dat(i_axi_r_pack    ),
        .i_cdc_buf_active(axi_o_rbusy),
        .o_cdc_buf_active(axi_i_rbusy),
        .o_clk  (i_clk  ),
        .o_rst_n(i_rst_n),
        .o_vld(i_axi_rvalid  ), 
        .o_rdy(i_axi_rready  ), 
        .o_dat(o_axi_r_pack) 
      );
       end
       else begin: r_async_fifo_gen
      e603_subsys_gnrl_cdc_fifo
      # (
        .DP(ASYNC_FIFO_DP),
        .DP_PTR_W (ASYNC_FIFO_DP_PTR_W),
        .DW  (AXI_R_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_r_cdc_fifo (
        .i_clk  (o_clk  ),
        .i_rst_n(o_rst_n),
        .i_vld(o_axi_rvalid), 
        .i_rdy(o_axi_rready), 
        .i_dat(i_axi_r_pack    ),
        .i_cdc_fifo_active(axi_o_rbusy),
        .o_cdc_fifo_active(axi_i_rbusy),
        .o_clk  (i_clk  ),
        .o_rst_n(i_rst_n),
        .o_vld(i_axi_rvalid  ), 
        .o_rdy(i_axi_rready  ), 
        .o_dat(o_axi_r_pack) 
      );
       end
      end
      else begin: r_sync_gen
    assign axi_o_rbusy = o_axi_rvalid;
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_R_BUF_PACK)
    ) u_axi_r_fifo(
    .i_clk_en(icb_clk_en),
    .i_vld(o_axi_rvalid), 
    .i_rdy(o_axi_rready), 
    .i_dat(i_axi_r_pack    ),
    .o_clk_en(axi_bus_clk_en),
    .o_vld(i_axi_rvalid  ), 
    .o_rdy(i_axi_rready  ), 
    .o_dat(o_axi_r_pack),
    .o_fifo_active(axi_i_rbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
      end
    endgenerate
  assign axi_buf_pipe_i_active = axi_i_arbusy | axi_i_rbusy;
  assign axi_buf_pipe_o_active = axi_o_arbusy | axi_o_rbusy;
endmodule
module  e603_subsys_gnrl_axi_buf_write # (
  parameter PAYLOAD_NORST = 0,
  parameter ASYNC = 0,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 0,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter AXLEN_W = 8,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           i_axi_awready,
  input                            i_axi_awvalid,
  input [ID_W-1:0]                 i_axi_awid,
  input [AW-1:0]                   i_axi_awaddr,
  input [AXLEN_W-1:0]                      i_axi_awlen,
  input [CMD_SIZE_W-1:0]                      i_axi_awsize,
  input [1:0]                      i_axi_awburst,
  input                            i_axi_awlock,
  input [3:0]                      i_axi_awcache,
  input [2:0]                      i_axi_awprot,
  input [USR_W-1:0]                i_axi_awuser, 
  output                           i_axi_wready,
  input                            i_axi_wvalid,
  input [DW-1:0]                   i_axi_wdata,
  input [MW-1:0]                   i_axi_wstrb,
  input                            i_axi_wlast,
  input                            i_axi_bready,
  output                           i_axi_bvalid,
  output [ID_W-1:0]                i_axi_bid,
  output [USR_W-1:0]               i_axi_buser,
  output [1:0]                     i_axi_bresp,
  input                            o_axi_awready,
  output                           o_axi_awvalid,
  output[ID_W-1:0]                 o_axi_awid,
  output[AW-1:0]                   o_axi_awaddr,
  output[AXLEN_W-1:0]                      o_axi_awlen,
  output[CMD_SIZE_W-1:0]                      o_axi_awsize,
  output[1:0]                      o_axi_awburst,
  output                           o_axi_awlock,
  output[3:0]                      o_axi_awcache,
  output[2:0]                      o_axi_awprot,
  output[USR_W-1:0]                o_axi_awuser, 
  input                            o_axi_wready,
  output                           o_axi_wvalid,
  output[DW-1:0]                   o_axi_wdata,
  output[MW-1:0]                   o_axi_wstrb,
  output                           o_axi_wlast,
  output                           o_axi_bready,
  input                            o_axi_bvalid,
  input  [USR_W-1:0]               o_axi_buser,
  input  [ID_W-1:0]                o_axi_bid,
  input  [1:0]                     o_axi_bresp,
  input                            axi_bus_clk_en,
  input                            icb_clk_en,
  output                           axi_buf_pipe_i_active,
  output                           axi_buf_pipe_o_active,
  input  i_clk,
  input  i_rst_n,
  input  o_clk,
  input  o_rst_n,
  input  clk,
  input  rst_n
  );
  wire i_axi_awready_raw;
  wire i_axi_awvalid_raw;
  wire i_axi_wready_raw;
  wire i_axi_wvalid_raw;
  assign i_axi_awvalid_raw = (~reset_flag_r) & i_axi_awvalid    ;
  assign i_axi_awready     = (~reset_flag_r) & i_axi_awready_raw;
  assign i_axi_wvalid_raw  = (~reset_flag_r) & i_axi_wvalid    ;
  assign i_axi_wready      = (~reset_flag_r) & i_axi_wready_raw;
    localparam AXI_AW_BUF_PACK = ID_W+AW+AXLEN_W+CMD_SIZE_W+2+1+3+4+USR_W;
    wire [AXI_AW_BUF_PACK-1:0] i_axi_aw_pack = {
                                             i_axi_awid    ,  
                                             i_axi_awaddr  ,
                                             i_axi_awlen   ,
                                             i_axi_awsize  ,
                                             i_axi_awburst ,
                                             i_axi_awlock  ,
                                             i_axi_awcache ,
                                             i_axi_awprot  ,
                                             i_axi_awuser   
                                            };
    wire [AXI_AW_BUF_PACK-1:0] o_axi_aw_pack ;
    assign  { 
              o_axi_awid    , 
              o_axi_awaddr  , 
              o_axi_awlen   , 
              o_axi_awsize  , 
              o_axi_awburst , 
              o_axi_awlock  , 
              o_axi_awcache , 
              o_axi_awprot  , 
              o_axi_awuser    
            } = o_axi_aw_pack ;
    wire axi_i_awbusy ; 
    wire axi_o_awbusy ; 
    generate 
      if(ASYNC == 1) begin: aw_async_gen
        if(ASYNC_FIFO == 0) begin: aw_async_buf_gen
      e603_subsys_gnrl_cdc_buf
      # (
        .DW  (AXI_AW_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_aw_cdc_buf (
        .i_clk  (i_clk  ),
        .i_rst_n(i_rst_n),
        .i_vld  (i_axi_awvalid_raw  ), 
        .i_rdy  (i_axi_awready_raw  ), 
        .i_dat  (i_axi_aw_pack),
        .i_cdc_buf_active(axi_i_awbusy),
        .o_cdc_buf_active(axi_o_awbusy),
        .o_clk  (o_clk  ),
        .o_rst_n(o_rst_n),
        .o_vld  (o_axi_awvalid), 
        .o_rdy  (o_axi_awready), 
        .o_dat  (o_axi_aw_pack) 
      );
       end
       else begin: aw_async_fifo_gen
      e603_subsys_gnrl_cdc_fifo
      # (
        .DP(ASYNC_FIFO_DP),
        .DP_PTR_W(ASYNC_FIFO_DP_PTR_W),
        .DW  (AXI_AW_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_aw_cdc_fifo (
        .i_clk  (i_clk  ),
        .i_rst_n(i_rst_n),
        .i_vld  (i_axi_awvalid_raw  ), 
        .i_rdy  (i_axi_awready_raw  ), 
        .i_dat  (i_axi_aw_pack),
        .i_cdc_fifo_active(axi_i_awbusy),
        .o_cdc_fifo_active(axi_o_awbusy),
        .o_clk  (o_clk  ),
        .o_rst_n(o_rst_n),
        .o_vld  (o_axi_awvalid), 
        .o_rdy  (o_axi_awready), 
        .o_dat  (o_axi_aw_pack) 
      );
       end
      end
      else begin: aw_sync_gen
     assign axi_i_awbusy = i_axi_awvalid_raw;
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_AW_BUF_PACK)
    ) u_axi_aw_fifo(
    .i_clk_en(axi_bus_clk_en), 
    .i_vld(i_axi_awvalid_raw  ), 
    .i_rdy(i_axi_awready_raw  ), 
    .i_dat(i_axi_aw_pack),
    .o_clk_en(icb_clk_en),
    .o_vld(o_axi_awvalid), 
    .o_rdy(o_axi_awready), 
    .o_dat(o_axi_aw_pack    ),
    .o_fifo_active(axi_o_awbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
      end
    endgenerate
    localparam AXI_W_BUF_PACK = DW+MW+1;
    wire [AXI_W_BUF_PACK-1:0] i_axi_w_pack = {
                                             i_axi_wdata      , 
                                             i_axi_wstrb      , 
                                             i_axi_wlast        
                                            };
    wire [AXI_W_BUF_PACK-1:0] o_axi_w_pack ;
    assign  { 
              o_axi_wdata  , 
              o_axi_wstrb  , 
              o_axi_wlast    
            } = o_axi_w_pack ;
    wire axi_i_wbusy ; 
    wire axi_o_wbusy ; 
    generate 
      if(ASYNC == 1) begin: w_async_gen
        if(ASYNC_FIFO == 0) begin: w_async_buf_gen
      e603_subsys_gnrl_cdc_buf
      # (
        .DW     (AXI_W_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_w_cdc_buf (
        .i_clk  (i_clk  ),
        .i_rst_n(i_rst_n),
        .i_vld  (i_axi_wvalid_raw  ), 
        .i_rdy  (i_axi_wready_raw  ), 
        .i_dat  (i_axi_w_pack),
        .i_cdc_buf_active(axi_i_wbusy),
        .o_cdc_buf_active(axi_o_wbusy),
        .o_clk  (o_clk  ),
        .o_rst_n(o_rst_n),
        .o_vld(o_axi_wvalid), 
        .o_rdy(o_axi_wready), 
        .o_dat(o_axi_w_pack    ) 
      );
       end
       else begin: w_async_fifo_gen
      e603_subsys_gnrl_cdc_fifo
      # (
        .DP(ASYNC_FIFO_DP),
        .DP_PTR_W(ASYNC_FIFO_DP_PTR_W),
        .DW     (AXI_W_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_w_cdc_fifo (
        .i_clk  (i_clk  ),
        .i_rst_n(i_rst_n),
        .i_vld  (i_axi_wvalid_raw  ), 
        .i_rdy  (i_axi_wready_raw  ), 
        .i_dat  (i_axi_w_pack),
        .i_cdc_fifo_active(axi_i_wbusy),
        .o_cdc_fifo_active(axi_o_wbusy),
        .o_clk  (o_clk  ),
        .o_rst_n(o_rst_n),
        .o_vld(o_axi_wvalid), 
        .o_rdy(o_axi_wready), 
        .o_dat(o_axi_w_pack    ) 
      );
       end
      end
      else begin: w_sync_gen
     assign axi_i_wbusy = i_axi_wvalid_raw;
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_W_BUF_PACK)
    ) u_axi_w_fifo(
    .i_clk_en(axi_bus_clk_en),
    .i_vld(i_axi_wvalid_raw  ), 
    .i_rdy(i_axi_wready_raw  ), 
    .i_dat(i_axi_w_pack),
    .o_clk_en(icb_clk_en),
    .o_vld(o_axi_wvalid), 
    .o_rdy(o_axi_wready), 
    .o_dat(o_axi_w_pack    ),
    .o_fifo_active(axi_o_wbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
      end
    endgenerate
    localparam AXI_B_BUF_PACK = USR_W + ID_W+2;
    wire [AXI_B_BUF_PACK-1:0] o_axi_b_pack = {
                                             o_axi_buser  ,  
                                             o_axi_bid  ,  
                                             o_axi_bresp        
                                            };
    wire [AXI_B_BUF_PACK-1:0] i_axi_b_pack ;
    assign  { 
              i_axi_buser    , 
              i_axi_bid    , 
              i_axi_bresp    
            } = i_axi_b_pack ;
    wire axi_i_bbusy ; 
    wire axi_o_bbusy ; 
    generate 
      if(ASYNC == 1) begin: b_async_gen
        if(ASYNC_FIFO == 0) begin: b_async_buf_gen
      e603_subsys_gnrl_cdc_buf
      # (
        .DW     (AXI_B_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_b_cdc_buf(
        .i_clk  (o_clk  ),
        .i_rst_n(o_rst_n),
        .i_vld  (o_axi_bvalid), 
        .i_rdy  (o_axi_bready), 
        .i_dat  (o_axi_b_pack    ),
        .i_cdc_buf_active(axi_o_bbusy),
        .o_cdc_buf_active(axi_i_bbusy),
        .o_clk  (i_clk  ),
        .o_rst_n(i_rst_n),
        .o_vld  (i_axi_bvalid  ), 
        .o_rdy  (i_axi_bready  ), 
        .o_dat  (i_axi_b_pack) 
      );
       end
       else begin: b_async_fifo_gen
      e603_subsys_gnrl_cdc_fifo
      # (
        .DP(ASYNC_FIFO_DP),
        .DP_PTR_W(ASYNC_FIFO_DP_PTR_W),
        .DW     (AXI_B_BUF_PACK),
        .SYNC_DP(SYNC_DP)
      ) u_axi_b_cdc_fifo(
        .i_clk  (o_clk  ),
        .i_rst_n(o_rst_n),
        .i_vld  (o_axi_bvalid), 
        .i_rdy  (o_axi_bready), 
        .i_dat  (o_axi_b_pack    ),
        .i_cdc_fifo_active(axi_o_bbusy),
        .o_cdc_fifo_active(axi_i_bbusy),
        .o_clk  (i_clk  ),
        .o_rst_n(i_rst_n),
        .o_vld  (i_axi_bvalid  ), 
        .o_rdy  (i_axi_bready  ), 
        .o_dat  (i_axi_b_pack) 
      );
       end
      end
      else begin: b_sync_gen
     assign axi_o_bbusy = o_axi_bvalid;
    e603_subsys_gnrl_ratio_fifo # (
        .PAYLOAD_NORST(PAYLOAD_NORST),
      .I_SUPPORT_RATIO (1),
      .O_SUPPORT_RATIO (1),
      .DP  (RATIO_FIFO_DP),
      .DW  (AXI_B_BUF_PACK)
    ) u_axi_b_fifo(
    .i_clk_en(icb_clk_en),
    .i_vld(o_axi_bvalid), 
    .i_rdy(o_axi_bready), 
    .i_dat(o_axi_b_pack    ),
    .o_clk_en(axi_bus_clk_en),
    .o_vld(i_axi_bvalid  ), 
    .o_rdy(i_axi_bready  ), 
    .o_dat(i_axi_b_pack),
    .o_fifo_active(axi_i_bbusy),
    .clk  (clk  ),
    .rst_n(rst_n)  
   );
      end
    endgenerate
   assign axi_buf_pipe_i_active = axi_i_awbusy | axi_i_wbusy | axi_i_bbusy;
   assign axi_buf_pipe_o_active = axi_o_awbusy | axi_o_wbusy | axi_o_bbusy;
endmodule
module  e603_subsys_gnrl_axi2ficb_write_async # (
  parameter ALLOW_FIX_BURST = 0,
  parameter SYNC_DP = 2,
  parameter ASYNC_FIFO = 0,
  parameter ASYNC_FIFO_DP = 0,
  parameter ASYNC_FIFO_DP_PTR_W = 0,
  parameter RATIO_FIFO_DP = 2,
  parameter CMD_SIZE_W = 3,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  input  reset_flag_r,
  output                           axi_awready,
  input                            axi_awvalid,
  input [ID_W-1:0]                 axi_awid,
  input [AW-1:0]                   axi_awaddr,
  input [7:0]                      axi_awlen,
  input [CMD_SIZE_W-1:0]                      axi_awsize,
  input [1:0]                      axi_awburst,
  input                            axi_awlock,
  input [3:0]                      axi_awcache,
  input [2:0]                      axi_awprot,
  input [USR_W-1:0]                axi_awuser, 
  output                           axi_wready,
  input                            axi_wvalid,
  input [DW-1:0]                   axi_wdata,
  input [MW-1:0]                   axi_wstrb,
  input                            axi_wlast,
  input                            axi_bready,
  output                           axi_bvalid,
  output [USR_W-1:0]               axi_buser,
  output [ID_W-1:0]                axi_bid,
  output [1:0]                     axi_bresp,
  output                           icb_wcmd_sel,
  output                           icb_wcmd_valid,
  input                            icb_wcmd_ready,
  output [AW-1:0]                  icb_wcmd_addr,
  output                           icb_wcmd_read, 
  output [DW-1:0]                  icb_wcmd_wdata,
  output [MW-1:0]                  icb_wcmd_wmask,
  output [1:0]                     icb_wcmd_beat,
  output                           icb_wcmd_lock,
  output                           icb_wcmd_excl,
  output [CMD_SIZE_W-1:0]         icb_wcmd_size,
  output [7:0]                     icb_wcmd_xlen,
  output [1:0]                     icb_wcmd_xburst,
  output [1:0]                     icb_wcmd_modes,
  output                           icb_wcmd_dmode,
  output [2:0]                     icb_wcmd_attri,
  output [USR_W-1:0]               icb_wcmd_usr,
  input                            icb_wrsp_valid,
  output                           icb_wrsp_ready,
  input                            icb_wrsp_err,
  input                            icb_wrsp_excl_ok,
  input [USR_W-1:0]                icb_wrsp_usr,
  output                           axi2icb_write_axi_active,
  output                           axi2icb_write_icb_active,
  input icb_clk  ,
  input icb_rst_n,  
  input async_axi_clk  ,
  input async_axi_rst_n  
  );
  wire                           o_axi_awready;
  wire                           o_axi_awvalid;
  wire[ID_W-1:0]                 o_axi_awid;
  wire[AW-1:0]                   o_axi_awaddr;
  wire[7:0]                      o_axi_awlen;
  wire[CMD_SIZE_W-1:0]                      o_axi_awsize;
  wire[1:0]                      o_axi_awburst;
  wire                           o_axi_awlock;
  wire[3:0]                      o_axi_awcache;
  wire[2:0]                      o_axi_awprot;
  wire[USR_W-1:0]                o_axi_awuser; 
  wire                           o_axi_wready;
  wire                           o_axi_wvalid;
  wire[DW-1:0]                   o_axi_wdata;
  wire[MW-1:0]                   o_axi_wstrb;
  wire                           o_axi_wlast;
  wire                           o_axi_bready;
  wire                           o_axi_bvalid;
  wire [USR_W-1:0]               o_axi_buser;
  wire [ID_W-1:0]                o_axi_bid;
  wire [1:0]                     o_axi_bresp;
  wire axi_buf_pipe_i_active;
  wire axi_buf_pipe_o_active;
  e603_subsys_gnrl_axi_buf_write # (
     .ASYNC (1),
     .SYNC_DP (SYNC_DP),
     .ASYNC_FIFO (ASYNC_FIFO),
     .ASYNC_FIFO_DP (ASYNC_FIFO_DP),
     .ASYNC_FIFO_DP_PTR_W (ASYNC_FIFO_DP_PTR_W),
     .RATIO_FIFO_DP(0),
  .CMD_SIZE_W(CMD_SIZE_W),
    .AW   (AW   ),
    .DW   (DW   ),
    .MW   (MW   ),
    .ID_W (ID_W ),
    .USR_W(USR_W) 
  ) u_axi_buf_write (
    .reset_flag_r(reset_flag_r),
    .i_axi_awready   (axi_awready   ),
    .i_axi_awvalid   (axi_awvalid   ),
    .i_axi_awid      (axi_awid      ),
    .i_axi_awaddr    (axi_awaddr    ),
    .i_axi_awlen     (axi_awlen     ),
    .i_axi_awsize    (axi_awsize    ),
    .i_axi_awburst   (axi_awburst   ),
    .i_axi_awlock    (axi_awlock    ),
    .i_axi_awcache   (axi_awcache   ),
    .i_axi_awprot    (axi_awprot    ),
    .i_axi_awuser    (axi_awuser    ), 
    .i_axi_wready    (axi_wready    ),
    .i_axi_wvalid    (axi_wvalid    ),
    .i_axi_wdata     (axi_wdata     ),
    .i_axi_wstrb     (axi_wstrb     ),
    .i_axi_wlast     (axi_wlast     ),
    .i_axi_bready    (axi_bready    ),
    .i_axi_bvalid    (axi_bvalid    ),
    .i_axi_buser     (axi_buser     ),
    .i_axi_bid       (axi_bid       ),
    .i_axi_bresp     (axi_bresp     ),
    .o_axi_awready   (o_axi_awready   ),
    .o_axi_awvalid   (o_axi_awvalid   ),
    .o_axi_awid      (o_axi_awid      ),
    .o_axi_awaddr    (o_axi_awaddr    ),
    .o_axi_awlen     (o_axi_awlen     ),
    .o_axi_awsize    (o_axi_awsize    ),
    .o_axi_awburst   (o_axi_awburst   ),
    .o_axi_awlock    (o_axi_awlock    ),
    .o_axi_awcache   (o_axi_awcache   ),
    .o_axi_awprot    (o_axi_awprot    ),
    .o_axi_awuser    (o_axi_awuser    ), 
    .o_axi_wready    (o_axi_wready    ),
    .o_axi_wvalid    (o_axi_wvalid    ),
    .o_axi_wdata     (o_axi_wdata     ),
    .o_axi_wstrb     (o_axi_wstrb     ),
    .o_axi_wlast     (o_axi_wlast     ),
    .o_axi_bready    (o_axi_bready    ),
    .o_axi_bvalid    (o_axi_bvalid    ),
    .o_axi_bid       (o_axi_bid       ),
    .o_axi_buser     (o_axi_buser     ),
    .o_axi_bresp     (o_axi_bresp     ),
    .axi_buf_pipe_i_active  (axi_buf_pipe_i_active),
    .axi_buf_pipe_o_active  (axi_buf_pipe_o_active),
    .i_clk                (async_axi_clk  ),
    .i_rst_n              (async_axi_rst_n),
    .o_clk                (icb_clk  ),
    .o_rst_n              (icb_rst_n),
    .axi_bus_clk_en       (1'b1),
    .icb_clk_en       (1'b1),
    .clk                  (1'b0),
    .rst_n                (1'b0)  
  );
  wire o_axi2icb_write_active;
  e603_subsys_gnrl_axi2ficb_write # (
  .ALLOW_FIX_BURST(ALLOW_FIX_BURST),
  .CMD_SIZE_W(CMD_SIZE_W),
  .AW(AW),
  .DW(DW),
  .MW(MW),
  .RATIO_FIFO_DP(0),
  .FIFO_OUTS_NUM(FIFO_OUTS_NUM),
  .ID_W (ID_W),
  .USR_W (USR_W)
  ) u_axi2icb_write (
    .reset_flag_r (1'b0),
    .axi_awready   (o_axi_awready   ),
    .axi_awvalid   (o_axi_awvalid   ),
    .axi_awid      (o_axi_awid      ),
    .axi_awaddr    (o_axi_awaddr    ),
    .axi_awlen     (o_axi_awlen     ),
    .axi_awsize    (o_axi_awsize    ),
    .axi_awburst   (o_axi_awburst   ),
    .axi_awlock    (o_axi_awlock    ),
    .axi_awcache   (o_axi_awcache   ),
    .axi_awprot    (o_axi_awprot    ),
    .axi_awuser    (o_axi_awuser    ), 
    .axi_wready    (o_axi_wready    ),
    .axi_wvalid    (o_axi_wvalid    ),
    .axi_wdata     (o_axi_wdata     ),
    .axi_wstrb     (o_axi_wstrb     ),
    .axi_wlast     (o_axi_wlast     ),
    .axi_bready    (o_axi_bready    ),
    .axi_bvalid    (o_axi_bvalid    ),
    .axi_bid       (o_axi_bid       ),
    .axi_buser     (o_axi_buser     ),
    .axi_bresp     (o_axi_bresp     ),
    .icb_wcmd_sel   (icb_wcmd_sel),
    .icb_wcmd_valid (icb_wcmd_valid ),
    .icb_wcmd_ready (icb_wcmd_ready ),
    .icb_wcmd_addr  (icb_wcmd_addr  ),
    .icb_wcmd_read  (icb_wcmd_read  ), 
    .icb_wcmd_wdata (icb_wcmd_wdata ),
    .icb_wcmd_wmask (icb_wcmd_wmask ),
    .icb_wcmd_beat  (icb_wcmd_beat  ),
    .icb_wcmd_lock  (icb_wcmd_lock  ),
    .icb_wcmd_excl  (icb_wcmd_excl  ),
    .icb_wcmd_size  (icb_wcmd_size  ),
    .icb_wcmd_xlen  (icb_wcmd_xlen    ),
    .icb_wcmd_xburst(icb_wcmd_xburst  ),
    .icb_wcmd_modes (icb_wcmd_modes   ),
    .icb_wcmd_dmode (icb_wcmd_dmode   ),
    .icb_wcmd_attri (icb_wcmd_attri   ),
    .icb_wcmd_usr   (icb_wcmd_usr ),
    .icb_wrsp_valid  (icb_wrsp_valid  ),
    .icb_wrsp_ready  (icb_wrsp_ready  ),
    .icb_wrsp_err    (icb_wrsp_err    ),
    .icb_wrsp_excl_ok(icb_wrsp_excl_ok),
    .icb_wrsp_usr     (icb_wrsp_usr),
    .axi_bus_clk_en  (1'b1),
    .icb_clk_en  (1'b1),
    .axi2icb_write_active  (o_axi2icb_write_active),
    .clk   (icb_clk  ),
    .rst_n (icb_rst_n)
  );
  assign axi2icb_write_axi_active = axi_buf_pipe_i_active;
  assign axi2icb_write_icb_active = axi_buf_pipe_o_active | o_axi2icb_write_active;
endmodule
`include "global.v"
module e603_subsys_gnrl_ficb_id_gen # (
  parameter OUTS_FIFO_DP = 8,
  parameter ID_W = 32 
) (
  input              i_icb_cmd_valid, 
  input              i_icb_cmd_ready, 
  input  [ID_W -1:0] i_icb_cmd_id,
  input  [2    -1:0] i_icb_cmd_xburst,
  input  [2    -1:0] i_icb_cmd_beat,
  input  [3    -1:0] i_icb_cmd_size,
  input  [8    -1:0] i_icb_cmd_xlen,
  output [2    -1:0] o_icb_cmd_beat,
  output [8    -1:0] o_icb_cmd_xlen,
  output             ficb_id_gen_ready,
  input              i_icb_rsp_valid, 
  input              i_icb_rsp_ready, 
  output [ID_W -1:0] i_icb_rsp_id,
  output             i_icb_rsp_last,
  input  clk,  
  input  rst_n
  );
  wire i_icb_cmd_fixed = (i_icb_cmd_xburst == 2'b00);
  assign o_icb_cmd_beat = i_icb_cmd_fixed ? 2'b0 : i_icb_cmd_beat;
  assign o_icb_cmd_xlen = i_icb_cmd_fixed ? 8'b0 : i_icb_cmd_xlen;
  wire i_icb_cmd_last = i_icb_cmd_beat[1] | (i_icb_cmd_xlen == 8'd0);
  wire i_icb_cmd_hsked = i_icb_cmd_valid & i_icb_cmd_ready;
  wire i_icb_rsp_hsked = i_icb_rsp_valid & i_icb_rsp_ready;
  wire rspid_fifo_o_vld;
     e603_subsys_gnrl_fifo # (
        .REG_OUT(0),
        .CUT_READY (1),
        .DP  (OUTS_FIFO_DP+1),
        .DW  (ID_W+1
               )
      ) u_e603_subsys_gnrl_rspid_fifo (
        .i_vld(i_icb_cmd_hsked),
        .i_rdy(ficb_id_gen_ready),
        .i_dat({i_icb_cmd_last,i_icb_cmd_id
               }),
        .o_vld(rspid_fifo_o_vld),
        .o_rdy(i_icb_rsp_hsked),
        .o_dat({i_icb_rsp_last,i_icb_rsp_id
               } ),
        .clk  (clk),
        .rst_n(rst_n)
      );
endmodule
`include "global.v"
module e603_subsys_gnrl_pipe_stage # (
  parameter CUT_READY = 0,
  parameter PAYLOAD_NORST = 0,
  parameter DP = 1,
  parameter DW = 32,
  parameter EW = DP == 0 ? 1 : ((DW-1)/64+1) + 1
) (
  input           i_vld,
  output          i_rdy,
  input  [DW-1:0] i_dat,
  output          o_vld,
  input           o_rdy,
  output [DW-1:0] o_dat,
  input           clk,
  input           rst_n
);
  genvar i;
  generate 
  if(DP == 0) begin: gen_dp_eq_0
      assign o_vld = i_vld;
      assign i_rdy = o_rdy;
      assign o_dat = i_dat;
  end
  else begin: gen_dp_gt_0
      wire vld_set;
      wire vld_clr;
      wire vld_ena;
      wire vld_r;
      wire vld_nxt;
      assign vld_set = i_vld & i_rdy;
      assign vld_clr = o_vld & o_rdy;
      assign vld_ena = vld_set | vld_clr;
      assign vld_nxt = vld_set | (~vld_clr);
e603_subsys_gnrl_dfflr #(1) vld_dfflr (vld_ena, vld_nxt, vld_r, clk, rst_n);// VPP_NO_REG_PARSE
    if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_dffl #(DW) dat_dffl (vld_set, i_dat, o_dat, clk, rst_n);// VPP_NO_REG_PARSE
    end
    else begin: rst_gen
e603_subsys_gnrl_dfflr #(DW) dat_dfflr (vld_set, i_dat, o_dat, clk, rst_n);// VPP_NO_REG_PARSE
    end
      assign o_vld = vld_r;
      if(CUT_READY == 1) begin:gen_cut_ready
          assign i_rdy = (~vld_r);
      end
      else begin:gen_no_cut_ready
          assign i_rdy = (~vld_r) | vld_clr;
      end
  end
  endgenerate
endmodule
module e603_subsys_gnrl_sync # (
  parameter DP = 2,
  parameter DW = 32,
  parameter [DW-1:0] RST_VAL = {DW{1'b0}}
) (
  input  [DW-1:0] din_a,
  output [DW-1:0] dout,
  input           rst_n,
  input           clk
);
`ifdef SYNTHESIS
 e603_gnrl_tech_sync #(
  .DP      (DP),
  .DW      (DW),
  .RST_VAL (RST_VAL)
) u_sync (
  .din_a (din_a  ),
  .dout  (dout   ),
  .rst_n (rst_n  ),
  .clk   (clk    )
);
`else
  wire [DW-1:0] sync_dat [DP-1:0];
  genvar i;
  generate
  for(i=0;i<DP;i=i+1) begin:gen_sync
    if(i==0) begin:gen_i_is_0
      e603_subsys_gnrl_cdc_dffrs #(DW, RST_VAL) sync_gnrl_cdc_dest_dffrs(din_a,         sync_dat[0], clk, rst_n);  // VPP_NO_REG_PARSE
    end
    else begin:gen_i_is_not_0
e603_subsys_gnrl_dffrs #(DW, RST_VAL) sync_dffrs(sync_dat[i-1], sync_dat[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
  end
  endgenerate
  assign dout = sync_dat[DP-1];
`endif
endmodule
module e603_subsys_gnrl_bus_sync (
  clk_s
  , rst_s_n
  , bus_s
  , clk_d
  , rst_d_n
  , bus_d
);
  parameter DW = 8;
  parameter DP = 2;
  input           clk_s;
  input           rst_s_n;
  input  [DW-1:0] bus_s;
  input           clk_d;
  input           rst_d_n;
  output [DW-1:0] bus_d;
  wire          lvl_s;
  wire [DW-1:0] bus_s_r;
  wire          lvl_d2s;
  wire          qlf_s;
  wire          lvl_d;
  wire [DW-1:0] bus_d_r;
  wire          lvl_s2d;
  wire          qlf_d;
  e603_subsys_gnrl_sync  #(
  .DW(1),
  .DP(DP))
  U_qlf_d2s_sync (
  .clk(clk_s),
  .rst_n(rst_s_n),
  .din_a(lvl_d),
  .dout(lvl_d2s)
  );
  assign qlf_s = lvl_s ^~ lvl_d2s;
  wire lvl_s_nxt;
  assign lvl_s_nxt = qlf_s ^ lvl_s;
e603_subsys_gnrl_dffr #(1) U_lvl_s_dffr (lvl_s_nxt, lvl_s, clk_s, rst_s_n);// VPP_NO_REG_PARSE
  wire [DW-1:0] bus_s_r_nxt;
  assign bus_s_r_nxt = qlf_s ? bus_s : bus_s_r;
  e603_subsys_gnrl_cdc_dffr #(DW) U_bus_s_r_gnrl_cdc_dest_dffr (bus_s_r_nxt, bus_s_r, clk_s, rst_s_n);  // VPP_NO_REG_PARSE
  e603_subsys_gnrl_sync  #(
  .DW(1),
  .DP(DP))
  U_qlf_s2d_sync (
  .clk(clk_d),
  .rst_n(rst_d_n),
  .din_a(lvl_s),
  .dout(lvl_s2d)
  );
  assign qlf_d = lvl_d ^ lvl_s2d;
  wire lvl_d_nxt;
  assign lvl_d_nxt = qlf_d ^ lvl_d;
e603_subsys_gnrl_dffr #(1) U_lvl_d_dffr (lvl_d_nxt, lvl_d, clk_d, rst_d_n);// VPP_NO_REG_PARSE
  wire [DW-1:0] bus_d_r_nxt;
  assign bus_d_r_nxt = qlf_d ? bus_s_r : bus_d_r;
  e603_subsys_gnrl_cdc_dffr #(DW) U_bus_d_r_gnrl_cdc_dest_dffr (bus_d_r_nxt, bus_d_r, clk_d, rst_d_n); // VPP_NO_REG_PARSE
  assign bus_d = bus_d_r;
endmodule
module e603_subsys_gnrl_rrobin_1cycle # (
    parameter ARBT_NUM = 4
)(
  output rrobin_active,
  output[ARBT_NUM-1:0] grt_vec,
  input [ARBT_NUM-1:0] req_vec,
  input arbt_ena,
  input clk,
  input rst_n
);
wire               req_cflt;
wire               indic_ena;
wire [ARBT_NUM-1:0] indic_nxt;
wire [ARBT_NUM-1:0] indic_r;
wire [ARBT_NUM-1:0] req_vec_ored;
wire [ARBT_NUM-1:0] req_vec_ored_sft1;
genvar i;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored
    assign req_vec_ored[i] = |req_vec[i:0];
  end
endgenerate
assign req_vec_ored_sft1 = {req_vec_ored[ARBT_NUM-2:0],1'b0};
wire [ARBT_NUM-1:0] req_vec_msked_ored_sft1;
assign req_vec_msked_ored_sft1= req_vec_ored_sft1 & req_vec;
wire req_vec_is_1hot = ~(|req_vec_msked_ored_sft1);
wire req_vec_not_zeros = (|req_vec);
wire req_vec_not_1hot  = ~req_vec_is_1hot;
assign req_cflt = req_vec_not_zeros & req_vec_not_1hot;
assign indic_ena  = req_cflt & arbt_ena;
e603_subsys_gnrl_dfflrs #(ARBT_NUM) indic_dfflr (indic_ena, indic_nxt, indic_r, clk, rst_n);// VPP_NO_REG_PARSE
wire [ARBT_NUM-1:0] req_vec_msked_1;
wire [ARBT_NUM-1:0] req_vec_msked_2;
wire [ARBT_NUM-1:0] ored_vec_msked_1;
wire [ARBT_NUM-1:0] vec_1hot_1;
wire [ARBT_NUM-1:0] grt_vec_1;
wire [ARBT_NUM-1:0] ored_vec_msked_2;
wire [ARBT_NUM-1:0] vec_1hot_2;
wire [ARBT_NUM-1:0] grt_vec_2;
wire [ARBT_NUM-1:0] req_vec_real;
assign rrobin_active = 1'b0;
assign req_vec_real = req_vec;
assign req_vec_msked_1 = indic_r & req_vec_real;
assign req_vec_msked_2 = (~indic_r) & req_vec_real;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored_vec_msked
    if(i==0) begin: gen_i_eq0
      assign ored_vec_msked_1[0] = req_vec_msked_1[0];
      assign ored_vec_msked_2[0] = req_vec_msked_2[0];
      assign vec_1hot_1[0] = ored_vec_msked_1[0];
      assign vec_1hot_2[0] = ored_vec_msked_2[0];
    end
    else begin: gen_i_neq0
      assign ored_vec_msked_1[i] = |req_vec_msked_1[i:0];
      assign ored_vec_msked_2[i] = |req_vec_msked_2[i:0];
      assign vec_1hot_1[i] = (~ored_vec_msked_1[i-1]) & ored_vec_msked_1[i];
      assign vec_1hot_2[i] = (~ored_vec_msked_2[i-1]) & ored_vec_msked_2[i];
    end
  end
endgenerate
assign grt_vec_1 = vec_1hot_1;
assign grt_vec_2 = vec_1hot_2;
wire grt_sel = |(indic_r & req_vec_real);
assign grt_vec = grt_sel ?  grt_vec_1 : grt_vec_2;
assign indic_nxt = grt_sel ?  {ored_vec_msked_1[ARBT_NUM-2:0],1'b0} : {ored_vec_msked_2[ARBT_NUM-2:0],1'b0};
endmodule
module e603_subsys_gnrl_rrobin_1cycle_da # (
    parameter ARBT_NUM = 4
)(
  output rrobin_active,
  output[ARBT_NUM-1:0] grt_vec,
  input [ARBT_NUM-1:0] req_vec,
  input [ARBT_NUM-1:0] buz_vec,
  input arbt_ena,
  input arbt_rply,
  input clk,
  input rst_n
);
wire                req_cflt;
wire [ARBT_NUM-1:0] req_vec_ored;
wire [ARBT_NUM-1:0] req_vec_ored_sft1;
genvar i;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored
    assign req_vec_ored[i] = |req_vec[i:0];
  end
endgenerate
assign req_vec_ored_sft1 = {req_vec_ored[ARBT_NUM-2:0],1'b0};
wire [ARBT_NUM-1:0] req_vec_msked_ored_sft1 = req_vec_ored_sft1 & req_vec;
wire req_vec_is_1hot = ~(|req_vec_msked_ored_sft1);
wire req_vec_not_zeros = (|req_vec);
wire req_vec_not_1hot  = ~req_vec_is_1hot;
assign req_cflt = req_vec_not_zeros & req_vec_not_1hot;
wire                indic_ena;
wire [ARBT_NUM-1:0] indic_nxt;
wire [ARBT_NUM-1:0] indic_r;
wire                indic_p_ena;
wire [ARBT_NUM-1:0] indic_p_nxt;
wire [ARBT_NUM-1:0] indic_p_r;
wire                indic_p1h_ena;
wire [ARBT_NUM-1:0] indic_p1h_nxt;
wire [ARBT_NUM-1:0] indic_p1h_r;
wire                indic_p1s_ena;
wire [ARBT_NUM-1:0] indic_p1s_nxt;
wire [ARBT_NUM-1:0] indic_p1s_r;
wire                indic_p1s_vld_r;
wire                indic_p1s_vld_nxt;
wire                indic_p1s_vld_ena;
wire                indic_p1s_rst_r;
wire                indic_p1s_rst_nxt;
wire                indic_p1s_rst_ena;
e603_subsys_gnrl_dfflrs #(ARBT_NUM) indic_dfflr (indic_ena, indic_nxt, indic_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflrs #(ARBT_NUM) indic_p_dfflr (indic_p_ena, indic_p_nxt, indic_p_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflrs #(ARBT_NUM, {{(ARBT_NUM-1){1'b0}}, 1'b1}) indic_p1h_dfflr (indic_p1h_ena, indic_p1h_nxt, indic_p1h_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflrs #(ARBT_NUM, {{(ARBT_NUM-1){1'b0}}, 1'b1}) indic_p1s_dfflr (indic_p1s_ena, indic_p1s_nxt, indic_p1s_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(1) indic_p1s_vld_dfflr (indic_p1s_vld_ena, indic_p1s_vld_nxt, indic_p1s_vld_r, clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr #(1) indic_p1s_rst_dfflr (indic_p1s_rst_ena, indic_p1s_rst_nxt, indic_p1s_rst_r, clk, rst_n);// VPP_NO_REG_PARSE
wire [ARBT_NUM-1:0] req_vec_msked_1;
wire [ARBT_NUM-1:0] req_vec_msked_2;
wire [ARBT_NUM-1:0] req_vec_msked_3;
wire [ARBT_NUM-1:0] req_vec_msked_4;
wire [ARBT_NUM-1:0] ored_vec_msked_1;
wire [ARBT_NUM-1:0] ored_vec_msked_2;
wire [ARBT_NUM-1:0] ored_vec_msked_3;
wire [ARBT_NUM-1:0] ored_vec_msked_4;
wire [ARBT_NUM-1:0] vec_1hot_1;
wire [ARBT_NUM-1:0] vec_1hot_2;
wire [ARBT_NUM-1:0] vec_1hot_3;
wire [ARBT_NUM-1:0] vec_1hot_4;
assign rrobin_active = 1'b0;
assign req_vec_msked_1 = indic_r & req_vec;
assign req_vec_msked_2 = (~indic_r) & req_vec;
assign req_vec_msked_3 = indic_p_r & buz_vec;
assign req_vec_msked_4 = (~indic_p_r) & buz_vec;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored_vec_msked
    if(i==0) begin: gen_i_eq0
      assign ored_vec_msked_1[0] = req_vec_msked_1[0];
      assign ored_vec_msked_2[0] = req_vec_msked_2[0];
      assign ored_vec_msked_3[0] = req_vec_msked_3[0];
      assign ored_vec_msked_4[0] = req_vec_msked_4[0];
      assign vec_1hot_1[0] = ored_vec_msked_1[0];
      assign vec_1hot_2[0] = ored_vec_msked_2[0];
      assign vec_1hot_3[0] = ored_vec_msked_3[0];
      assign vec_1hot_4[0] = ored_vec_msked_4[0];
    end
    else begin: gen_i_neq0
      assign ored_vec_msked_1[i] = |req_vec_msked_1[i:0];
      assign ored_vec_msked_2[i] = |req_vec_msked_2[i:0];
      assign ored_vec_msked_3[i] = |req_vec_msked_3[i:0];
      assign ored_vec_msked_4[i] = |req_vec_msked_4[i:0];
      assign vec_1hot_1[i] = (~ored_vec_msked_1[i-1]) & ored_vec_msked_1[i];
      assign vec_1hot_2[i] = (~ored_vec_msked_2[i-1]) & ored_vec_msked_2[i];
      assign vec_1hot_3[i] = (~ored_vec_msked_3[i-1]) & ored_vec_msked_3[i];
      assign vec_1hot_4[i] = (~ored_vec_msked_4[i-1]) & ored_vec_msked_4[i];
    end
  end
endgenerate
wire grt_sel1 = |req_vec_msked_1;
wire grt_sel3 = |req_vec_msked_3;
wire grt_sel4 = |(req_vec & indic_p1h_r);
wire [ARBT_NUM-1:0] grt_vec_np = grt_sel1 ? vec_1hot_1: vec_1hot_2;
wire grt_np_is_p = |(indic_p1h_r & grt_vec_np);
wire p_deasserted = ~(|(indic_p1h_r & buz_vec));
assign grt_vec = grt_sel4 ? indic_p1h_r : grt_vec_np;
wire [ARBT_NUM-1:0] ored_vec_msked_sel = grt_sel1 ? ored_vec_msked_1 : ored_vec_msked_2;
assign indic_ena = (~grt_sel4 | grt_np_is_p) & req_cflt & arbt_ena;
assign indic_nxt = {ored_vec_msked_sel[ARBT_NUM-2:0],1'b0};
wire [ARBT_NUM-1:0] ored_vec_msked_pri = grt_sel3 ? ored_vec_msked_3 : ored_vec_msked_4;
wire [ARBT_NUM-1:0] ored_vec_msked_pri_1h = grt_sel3 ? vec_1hot_3 : vec_1hot_4;
wire   indic_p_pass = grt_sel4 & arbt_ena;
wire   indic_p_rply = indic_p1s_vld_r & arbt_rply;
wire   indic_p_rstr = indic_p1s_rst_r & indic_p_pass;
wire   indic_p_rr   = indic_p_rply | indic_p_rstr;
assign indic_p_ena = ((grt_sel4 & ~indic_p_rr) | p_deasserted) & arbt_ena;
assign indic_p_nxt = {ored_vec_msked_pri[ARBT_NUM-2:0],1'b0};
assign indic_p1h_ena = indic_p_ena | indic_p_rr;
assign indic_p1h_nxt = indic_p_rr ? indic_p1s_r : ored_vec_msked_pri_1h;
assign indic_p1s_ena = indic_p_pass | indic_p_rply;
assign indic_p1s_nxt = indic_p1h_r;
assign indic_p1s_vld_ena = arbt_ena & req_vec_not_zeros;
assign indic_p1s_vld_nxt = grt_sel4;
assign indic_p1s_rst_ena = indic_p_rr;
assign indic_p1s_rst_nxt = indic_p_rply;
endmodule
module e603_subsys_gnrl_rrobin # (
    parameter ARBT_NUM = 4
)(
  output rrobin_active,
  output[ARBT_NUM-1:0] grt_vec,
  input [ARBT_NUM-1:0] req_vec,
  input arbt_ena,
  input clk,
  input rst_n
);
wire               req_cflt;
wire               indic_ena;
wire               indic_ovf;
wire [ARBT_NUM-1:0] indic_nxt;
wire [ARBT_NUM-1:0] indic_r;
wire [ARBT_NUM-1:0] req_vec_ored;
wire [ARBT_NUM-1:0] req_vec_ored_sft1;
genvar i;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored
    assign req_vec_ored[i] = |req_vec[i:0];
  end
endgenerate
assign req_vec_ored_sft1 = {req_vec_ored[ARBT_NUM-2:0],1'b0};
wire [ARBT_NUM-1:0] req_vec_msked_ored_sft1;
assign req_vec_msked_ored_sft1= req_vec_ored_sft1 & req_vec;
wire req_vec_is_1hot = ~(|req_vec_msked_ored_sft1);
wire req_vec_not_zeros = (|req_vec);
wire req_vec_not_1hot  = ~req_vec_is_1hot;
assign req_cflt = req_vec_not_zeros & req_vec_not_1hot;
assign indic_ena  = req_cflt & arbt_ena;
generate
  if(ARBT_NUM == 2) begin: gen_arbtnum_eq_2
    assign indic_ovf = ~(indic_r[0]);
  end
  else begin: gen_arbtnum_ueq_2
    assign indic_ovf = ~(|indic_r[ARBT_NUM-2:0]);
  end
endgenerate
e603_subsys_gnrl_dfflrs #(ARBT_NUM) indic_dfflr (indic_ena, indic_nxt, indic_r, clk, rst_n);// VPP_NO_REG_PARSE
wire [ARBT_NUM-1:0] req_vec_msked_1;
wire [ARBT_NUM-1:0] req_vec_msked_2;
wire [ARBT_NUM-1:0] ored_vec_msked_1;
wire [ARBT_NUM-1:0] vec_1hot_1;
wire [ARBT_NUM-1:0] grt_vec_1;
wire [ARBT_NUM-1:0] ored_vec_msked_2;
wire [ARBT_NUM-1:0] vec_1hot_2;
wire [ARBT_NUM-1:0] grt_vec_2;
wire [ARBT_NUM-1:0] mask_r;
wire [ARBT_NUM-1:0] mask_nxt;
wire mask_ena;
wire mask_set;
wire mask_clr;
wire [ARBT_NUM-1:0] req_vec_real;
assign mask_set = (|grt_vec) & (~arbt_ena);
assign mask_clr = (arbt_ena | (~(|req_vec_real))) & (|mask_r);
assign mask_ena = mask_set | mask_clr;
assign mask_nxt = mask_clr ? {ARBT_NUM{1'b0}} : (~grt_vec);
e603_subsys_gnrl_dfflr #(ARBT_NUM) mask_dfflr (mask_ena, mask_nxt, mask_r, clk, rst_n);// VPP_NO_REG_PARSE
assign rrobin_active = (|mask_r);
assign req_vec_real = req_vec & (~mask_r);
assign req_vec_msked_1 = indic_r & req_vec_real;
assign req_vec_msked_2 = (~indic_r) & req_vec_real;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored_vec_msked
    if(i==0) begin: gen_i_eq0
      assign ored_vec_msked_1[0] = req_vec_msked_1[0];
      assign ored_vec_msked_2[0] = req_vec_msked_2[0];
      assign vec_1hot_1[0] = ored_vec_msked_1[0];
      assign vec_1hot_2[0] = ored_vec_msked_2[0];
    end
    else begin: gen_i_neq0
      assign ored_vec_msked_1[i] = |req_vec_msked_1[i:0];
      assign ored_vec_msked_2[i] = |req_vec_msked_2[i:0];
      assign vec_1hot_1[i] = (~ored_vec_msked_1[i-1]) & ored_vec_msked_1[i];
      assign vec_1hot_2[i] = (~ored_vec_msked_2[i-1]) & ored_vec_msked_2[i];
    end
  end
endgenerate
assign grt_vec_1 = vec_1hot_1;
assign grt_vec_2 = vec_1hot_2;
wire grt_sel = |(indic_r & req_vec_real);
assign grt_vec = grt_sel ?  grt_vec_1 : grt_vec_2;
assign indic_nxt = grt_sel ?  {ored_vec_msked_1[ARBT_NUM-2:0],1'b0} : {ored_vec_msked_2[ARBT_NUM-2:0],1'b0};
endmodule
module e603_subsys_gnrl_rrobin_cut # (
    parameter ARBT_NUM = 4
)(
  output rrobin_active,
  output[ARBT_NUM-1:0] grt_vec,
  input [ARBT_NUM-1:0] req_vec,
  input arbt_ena,
  input [ARBT_NUM-1:0] req_mask,
  input req_mask_set,
  input clk,
  input rst_n
);
  wire req_mask_ored = (|req_mask);
  wire req_mask_set_real = req_mask_set & (~req_mask_ored);
wire [ARBT_NUM-1:0] grt_vec_old;
wire               req_cflt;
wire               indic_ena;
wire               indic_ovf;
wire [ARBT_NUM-1:0] indic_nxt;
wire [ARBT_NUM-1:0] indic_r;
wire [ARBT_NUM-1:0] req_vec_ored;
wire [ARBT_NUM-1:0] req_vec_ored_sft1;
genvar i;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored
    assign req_vec_ored[i] = |req_vec[i:0];
  end
endgenerate
assign req_vec_ored_sft1 = {req_vec_ored[ARBT_NUM-2:0],1'b0};
wire [ARBT_NUM-1:0] req_vec_msked_ored_sft1;
assign req_vec_msked_ored_sft1= req_vec_ored_sft1 & req_vec;
wire req_vec_is_1hot = ~(|req_vec_msked_ored_sft1);
wire req_vec_not_zeros = (|req_vec);
wire req_vec_not_1hot  = ~req_vec_is_1hot;
assign req_cflt = req_vec_not_zeros & req_vec_not_1hot;
wire empty_grt;
assign indic_ena  = (req_cflt & arbt_ena) | empty_grt;
generate
  if(ARBT_NUM == 2) begin: gen_arbtnum_eq_2
    assign indic_ovf = ~(indic_r[0]);
  end
  else begin: gen_arbtnum_ueq_2
    assign indic_ovf = ~(|indic_r[ARBT_NUM-2:0]);
  end
endgenerate
wire [ARBT_NUM-1:0] indic_r_1hot;
e603_subsys_gnrl_dfflrs #(ARBT_NUM) indic_dfflr (indic_ena, indic_nxt, indic_r, clk, rst_n);// VPP_NO_REG_PARSE
wire [ARBT_NUM-1:0] req_vec_msked_1;
wire [ARBT_NUM-1:0] req_vec_msked_2;
wire [ARBT_NUM-1:0] ored_vec_msked_1;
wire [ARBT_NUM-1:0] vec_1hot_1;
wire [ARBT_NUM-1:0] ored_vec_msked_2;
wire [ARBT_NUM-1:0] vec_1hot_2;
wire [ARBT_NUM-1:0] grt_vec_1;
wire [ARBT_NUM-1:0] grt_vec_2;
wire [ARBT_NUM-1:0] req_hck_msked_1;
wire [ARBT_NUM-1:0] req_hck_msked_2;
wire [ARBT_NUM-1:0] ored_hck_msked_1;
wire [ARBT_NUM-1:0] hck_1hot_1;
wire [ARBT_NUM-1:0] ored_hck_msked_2;
wire [ARBT_NUM-1:0] hck_1hot_2;
wire [ARBT_NUM-1:0] mask_r;
wire [ARBT_NUM-1:0] mask_nxt;
wire mask_ena;
wire mask_set;
wire mask_clr;
wire [ARBT_NUM-1:0] req_vec_real;
wire [ARBT_NUM-1:0] req_hck_real;
wire [ARBT_NUM-1:0] req_vec_masked;
assign req_vec_masked = req_vec & mask_r;
assign mask_set = (|grt_vec_old) & (~arbt_ena) & (~req_mask_ored);
assign mask_clr = (arbt_ena | (~(|req_vec_masked))) & (|mask_r);
assign mask_ena = mask_set | mask_clr;
assign mask_nxt = mask_clr ? {ARBT_NUM{1'b0}} : (~grt_vec_old);
e603_subsys_gnrl_dfflr #(ARBT_NUM) mask_dfflr (mask_ena, mask_nxt, mask_r, clk, rst_n);// VPP_NO_REG_PARSE
assign rrobin_active = (|mask_r);
wire mask_r_ored = rrobin_active;
assign req_vec_real = req_vec;
assign req_hck_real = req_vec_real & (~grt_vec);
assign req_vec_msked_1 = indic_r & req_vec_real;
assign req_vec_msked_2 = (~indic_r) & req_vec_real;
assign req_hck_msked_1 = indic_r & req_hck_real;
assign req_hck_msked_2 = (~indic_r) & req_hck_real;
generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:gen_ored_vec_msked
    if(i==0) begin: gen_i_eq0
      assign ored_vec_msked_1[0] = req_vec_msked_1[0];
      assign ored_vec_msked_2[0] = req_vec_msked_2[0];
      assign vec_1hot_1[0] = ored_vec_msked_1[0];
      assign vec_1hot_2[0] = ored_vec_msked_2[0];
      assign ored_hck_msked_1[0] = req_hck_msked_1[0];
      assign ored_hck_msked_2[0] = req_hck_msked_2[0];
      assign hck_1hot_1[0] = ored_hck_msked_1[0];
      assign hck_1hot_2[0] = ored_hck_msked_2[0];
      assign indic_r_1hot[0] = indic_r[0];
    end
    else begin: gen_i_neq0
      assign ored_vec_msked_1[i] = |req_vec_msked_1[i:0];
      assign ored_vec_msked_2[i] = |req_vec_msked_2[i:0];
      assign vec_1hot_1[i] = (~ored_vec_msked_1[i-1]) & ored_vec_msked_1[i];
      assign vec_1hot_2[i] = (~ored_vec_msked_2[i-1]) & ored_vec_msked_2[i];
      assign ored_hck_msked_1[i] = |req_hck_msked_1[i:0];
      assign ored_hck_msked_2[i] = |req_hck_msked_2[i:0];
      assign hck_1hot_1[i] = (~ored_hck_msked_1[i-1]) & ored_hck_msked_1[i];
      assign hck_1hot_2[i] = (~ored_hck_msked_2[i-1]) & ored_hck_msked_2[i];
      assign indic_r_1hot[i] = (~indic_r[i-1]) & indic_r[i];
    end
  end
endgenerate
wire grt_sel = |(indic_r & req_vec_real);
wire hck_sel = |(indic_r & req_hck_real);
assign grt_vec_1 = vec_1hot_1;
assign grt_vec_2 = vec_1hot_2;
    assign grt_vec = mask_r_ored ? (~mask_r) : req_mask_ored ? (~req_mask) : indic_r_1hot;
    assign grt_vec_old = grt_sel ?  grt_vec_1 : grt_vec_2;
    assign empty_grt = ((~(|(grt_vec & req_vec_real))) & (|req_vec_real)) 
                     & (~req_mask_ored) 
                     & (~mask_r_ored);
    assign indic_nxt = empty_grt ? (grt_sel ? {ored_vec_msked_1[ARBT_NUM-1:0]} : {ored_vec_msked_2[ARBT_NUM-1:0]}) :
                                   (hck_sel ? {ored_hck_msked_1[ARBT_NUM-1:0]} : {ored_hck_msked_2[ARBT_NUM-1:0]}) ;
endmodule
module e603_subsys_gnrl_rrobin_time # (
    parameter ARBT_NUM = 4
)(
  output rrobin_active,
  output[ARBT_NUM-1:0] grt_vec,
  input [ARBT_NUM-1:0] req_vec,
  input [ARBT_NUM-1:0] req_mask,
  input arbt_ena,
  input clk,
  input rst_n
);
  genvar i;
  wire [ARBT_NUM-1:0] i_grt_vec;
  wire [ARBT_NUM-1:0] i_req_vec;
  wire i_rrobin_active;
  wire req_mask_ored = (|req_mask);
  wire arbt_ena_msked = arbt_ena & req_mask_ored;
  e603_subsys_gnrl_rrobin # (
      .ARBT_NUM(ARBT_NUM)
  )u_gnrl_rrobin(
    .rrobin_active(i_rrobin_active),
    .grt_vec (i_grt_vec),
    .req_vec (i_req_vec),
    .arbt_ena(arbt_ena_msked),
    .clk     (clk     ),
    .rst_n   (rst_n   )
  );
  wire fifo_i_push;
  wire fifo_o_vld;
  wire fifo_o_pop;
  wire [ARBT_NUM-1:0] fifo_i_req_vec;
  wire [ARBT_NUM-1:0] fifo_o_req_vec;
  e603_subsys_gnrl_fifo # (
       .DP(ARBT_NUM+1),
       .DW(ARBT_NUM),
       .CUT_READY(1)
  ) u_arbt_pend_fifo(
    .i_vld   (fifo_i_push),
    .i_rdy   (),
    .i_dat   (fifo_i_req_vec),
    .o_vld   (fifo_o_vld),
    .o_rdy   (fifo_o_pop),
    .o_dat   (fifo_o_req_vec),
    .clk     (clk  ),
    .rst_n   (rst_n)
  );
  wire [ARBT_NUM-1:0] req_pend_r;
  wire [ARBT_NUM-1:0] req_pend_nxt;
  wire [ARBT_NUM-1:0] req_pend_ena;
  wire [ARBT_NUM-1:0] req_pend_set;
  wire [ARBT_NUM-1:0] req_pend_clr;
  wire [ARBT_NUM-1:0] req_pend_clr_raw;
  generate
    for(i = 0; i < ARBT_NUM; i = i+1)
    begin:gen_req_pend
        assign req_pend_set[i] = (~req_pend_r[i]) & (~(grt_vec[i] & arbt_ena)) & req_vec[i]
                               & (~(
                                    req_mask_ored ? grt_vec[i] : 1'b0
                                    )
                                 )
                               ;
        assign req_pend_clr_raw[i] = fifo_o_vld & fifo_o_req_vec[i] & ((grt_vec[i] & arbt_ena) | (~req_vec[i]));
        assign req_pend_clr[i] = req_pend_r[i] & req_pend_clr_raw[i];
        assign req_pend_ena[i] = req_pend_set[i] | req_pend_clr[i];
        assign req_pend_nxt[i] = (~req_pend_clr[i]);
e603_subsys_gnrl_dfflr #(1) req_pend_dfflr (req_pend_ena[i], req_pend_nxt[i], req_pend_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
  endgenerate
  assign fifo_i_push = (|req_pend_set);
  assign fifo_i_req_vec = req_pend_set;
  wire [ARBT_NUM-1:0] fifo_o_grted_vec_r;
  wire [ARBT_NUM-1:0] fifo_o_req_vec_real = req_vec & fifo_o_req_vec & (~fifo_o_grted_vec_r);
  assign fifo_o_pop = fifo_o_vld & (~(|fifo_o_req_vec_real));
  wire [ARBT_NUM-1:0] fifo_o_grted_vec_nxt;
  wire [ARBT_NUM-1:0] fifo_o_grted_vec_ena;
  wire [ARBT_NUM-1:0] fifo_o_grted_vec_set;
  wire [ARBT_NUM-1:0] fifo_o_grted_vec_clr;
  generate
    for(i = 0; i < ARBT_NUM; i = i+1)
    begin:gen_fifo_o_grted_vec
        assign fifo_o_grted_vec_set[i] = (~fifo_o_grted_vec_r[i]) & req_pend_clr_raw[i] & (~fifo_o_pop);
        assign fifo_o_grted_vec_clr[i] = fifo_o_grted_vec_r[i] & fifo_o_pop;
        assign fifo_o_grted_vec_ena[i] = fifo_o_grted_vec_set[i] | fifo_o_grted_vec_clr[i];
        assign fifo_o_grted_vec_nxt[i] = (~fifo_o_grted_vec_clr[i]);
e603_subsys_gnrl_dfflr #(1) fifo_o_grted_vec_dfflr (fifo_o_grted_vec_ena[i], fifo_o_grted_vec_nxt[i], fifo_o_grted_vec_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
  endgenerate
  assign i_req_vec =
      req_mask_ored ? {ARBT_NUM{1'b0}} :
      fifo_o_vld    ? fifo_o_req_vec_real :
                      req_vec;
  assign grt_vec = req_mask_ored ? (~req_mask) : i_grt_vec;
  assign rrobin_active = i_rrobin_active | fifo_o_vld;
endmodule
module e603_subsys_gnrl_cdc_tx
# (
  parameter PAYLOAD_NORST = 0,
  parameter DW = 32,
  parameter SYNC_DP = 2
) (
  input  i_vld,
  output i_rdy,
  input  [DW-1:0] i_dat,
  output o_vld,
  input  o_rdy_a,
  output [DW-1:0] o_dat,
  input  clk,
  input  rst_n
);
wire o_rdy_sync;
e603_subsys_gnrl_sync #(
    .DP(SYNC_DP),
    .DW(1)
) u_o_rdy_sync (
         .clk   (clk),
         .rst_n (rst_n),
         .din_a (o_rdy_a),
         .dout  (o_rdy_sync)
        );
wire vld_r;
wire [DW-1:0] dat_r;
wire vld_set = i_vld & i_rdy;
wire vld_clr = o_vld & o_rdy_sync;
wire vld_ena = vld_set | vld_clr;
wire vld_nxt = vld_set | (~vld_clr);
e603_subsys_gnrl_cdc_dfflr #(1) vld_dfflr(vld_ena, vld_nxt, vld_r, clk, rst_n); // VPP_NO_REG_PARSE
generate
if(PAYLOAD_NORST == 1) begin: no_rst_gen
e603_subsys_gnrl_cdc_dfflr #(DW) dat_dfflr(vld_set, i_dat, dat_r, clk, rst_n);  // VPP_NO_REG_PARSE
end
else begin: rst_gen
e603_subsys_gnrl_cdc_dffl #(DW) dat_dffl(vld_set, i_dat, dat_r, clk, rst_n);  // VPP_NO_REG_PARSE
end
endgenerate
wire o_rdy_sync_r;
e603_subsys_gnrl_dffr #(1) o_rdy_sync_dffr(o_rdy_sync, o_rdy_sync_r, clk, rst_n);// VPP_NO_REG_PARSE
wire o_rdy_nedge = (~o_rdy_sync) & o_rdy_sync_r;
wire nrdy_r;
wire nrdy_set = vld_set;
wire nrdy_clr = o_rdy_nedge;
wire nrdy_ena = nrdy_set | nrdy_clr;
wire nrdy_nxt = nrdy_set | (~nrdy_clr);
e603_subsys_gnrl_dfflr #(1) buf_nrdy_dfflr(nrdy_ena, nrdy_nxt, nrdy_r, clk, rst_n);// VPP_NO_REG_PARSE
assign o_vld = vld_r;
assign o_dat = dat_r;
assign i_rdy = (~nrdy_r) | nrdy_clr;
endmodule
module e603_subsys_gnrl_cdc_req_channel
# (
  parameter SYNC_DP = 2
) (
  input  req_i, 
  output req_o, 
  input  ack_a, 
  input  clk,
  input  rst_n 
);
  e603_subsys_gnrl_cdc_tx # (
     .DW      (1),
     .SYNC_DP (SYNC_DP)
   ) u_cdc_req_channel (
  .i_vld   (req_i),
  .i_rdy   (),
  .i_dat   (1'b0),
  .o_vld   (req_o),
  .o_rdy_a (ack_a),
  .o_dat   (),
  .clk     (clk),
  .rst_n   (rst_n)
);
endmodule
module e603_subsys_gnrl_bypbuf # (
  parameter PAYLOAD_NORST = 0,
  parameter DP = 1,
  parameter DW = 32
) (
  input           i_vld,
  output          i_rdy,
  input  [DW-1:0] i_dat,
  output          o_vld,
  input           o_rdy,
  output [DW-1:0] o_dat,
  output          fifo_o_vld,
  input           clk,
  input           rst_n
);
  wire          fifo_i_vld;
  wire          fifo_i_rdy;
  wire [DW-1:0] fifo_i_dat;
  wire          fifo_o_rdy;
  wire [DW-1:0] fifo_o_dat;
  e603_subsys_gnrl_fifo # (
       .PAYLOAD_NORST(PAYLOAD_NORST),
       .DP(DP),
       .DW(DW),
       .CUT_READY(1)
  ) u_bypbuf_fifo(
    .i_vld   (fifo_i_vld),
    .i_rdy   (fifo_i_rdy),
    .i_dat   (fifo_i_dat),
    .o_vld   (fifo_o_vld),
    .o_rdy   (fifo_o_rdy),
    .o_dat   (fifo_o_dat),
    .clk     (clk  ),
    .rst_n   (rst_n)
  );
  assign i_rdy = fifo_i_rdy;
  wire byp = i_vld & o_rdy & (~fifo_o_vld);
  assign fifo_o_rdy = o_rdy;
  assign o_vld = fifo_o_vld | i_vld;
  assign o_dat = fifo_o_vld ? fifo_o_dat : i_dat;
  assign fifo_i_dat  = i_dat;
  assign fifo_i_vld = i_vld & (~byp);
endmodule
module e603_subsys_gnrl_ratio_bypbuf # (
  parameter PAYLOAD_NORST = 0,
  parameter DP = 8,
  parameter DW = 32
) (
  input           clk_en,
  input           i_vld,
  output          i_rdy,
  input  [DW-1:0] i_dat,
  output          o_vld,
  input           o_rdy,
  output [DW-1:0] o_dat,
  input           clk,
  input           rst_n
);
  wire          fifo_i_vld;
  wire          fifo_i_rdy;
  wire [DW-1:0] fifo_i_dat;
  wire          fifo_o_vld;
  wire          fifo_o_rdy;
  wire [DW-1:0] fifo_o_dat;
  e603_subsys_gnrl_ratio_fifo # (
       .PAYLOAD_NORST(PAYLOAD_NORST),
       .I_SUPPORT_RATIO(1),
       .O_SUPPORT_RATIO(1),
       .DP(DP),
       .DW(DW)
  ) u_bypbuf_ratio_fifo(
    .i_clk_en(clk_en),
    .o_clk_en(clk_en),
    .i_vld   (fifo_i_vld),
    .i_rdy   (fifo_i_rdy),
    .i_dat   (fifo_i_dat),
    .o_vld   (fifo_o_vld),
    .o_rdy   (fifo_o_rdy),
    .o_dat   (fifo_o_dat),
    .o_fifo_active(),
    .clk     (clk  ),
    .rst_n   (rst_n)
  );
  assign i_rdy = fifo_i_rdy;
  wire byp = i_vld & o_rdy & (~fifo_o_vld);
  assign fifo_o_rdy = o_rdy;
  assign o_vld = fifo_o_vld | i_vld;
  assign o_dat = fifo_o_vld ? fifo_o_dat : i_dat;
  assign fifo_i_dat  = i_dat;
  assign fifo_i_vld = i_vld & (~byp);
endmodule
module e603_subsys_gnrl_stck # (
  parameter PAYLOAD_NORST = 0,
  parameter DP   = 8,
  parameter DW   = 32
) (
  input           i_wen,
  input  [DW-1:0] i_dat,
  input           o_ren,
  output [DW-1:0] o_dat,
  input           clk,
  input           rst_n
);
  wire [DW-1:0] stck_rf_r [DP-1:0];
  wire [DP-1:0] stck_rf_en;
  wire [DP:0] i_vec;
  wire [DP:0] o_vec;
  wire [DP:0] vec_nxt;
  wire [DP:0] vec_r;
  wire vec_en = (o_ren ^ i_wen );
  assign vec_nxt = i_wen ? (vec_r << 1) : (vec_r >> 1);
e603_subsys_gnrl_dfflrs #(1)  vec_0_dfflrs(vec_en, vec_nxt[0]   , vec_r[0]   , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP) vec_dp_dfflr(vec_en, vec_nxt[DP:1], vec_r[DP:1], clk, rst_n);// VPP_NO_REG_PARSE
  assign i_vec = vec_r; 
  assign o_vec = (vec_r >> 1); 
  genvar i;
  generate 
    for (i=0; i<DP; i=i+1) begin:gen_stck_rf
      assign stck_rf_en[i] = i_wen & i_vec[i];      
    if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_dffl  #(DW) stck_rf_dffl (stck_rf_en[i], i_dat, stck_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
    else begin: rst_gen
e603_subsys_gnrl_dfflr #(DW) stck_rf_dfflr(stck_rf_en[i], i_dat, stck_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
    end
  endgenerate
  integer j;
  reg [DW-1:0] mux_rdat;
  always @*
  begin : rd_port_PROC
    mux_rdat = {DW{1'b0}};
    for(j=0; j<DP; j=j+1) begin
      mux_rdat = mux_rdat | ({DW{o_vec[j]}} & stck_rf_r[j]);
    end
  end
  assign o_dat = mux_rdat;
endmodule
module e603_subsys_gnrl_ratio_fifo # (
  parameter PAYLOAD_NORST = 0,
  parameter I_SUPPORT_RATIO = 0,
  parameter O_SUPPORT_RATIO = 0,
  parameter REG_OUT = 0,
  parameter DP   = 8,
  parameter DW   = 32
) (
  input           i_clk_en,
  input           i_vld,
  output          i_rdy,
  input  [DW-1:0] i_dat,
  input           o_clk_en,
  output          o_vld,
  input           o_rdy,
  output [DW-1:0] o_dat,
  output          o_fifo_active,
  input           clk,
  input           rst_n
);
genvar i;
generate
  if(DP == 0) begin: gen_dp_eq1
     assign o_vld = i_vld;
     assign i_rdy = o_rdy;
     assign o_dat = i_dat;
     assign o_fifo_active =  i_vld;
  end
  else begin: gen_dp_gt0
    wire [DW-1:0] fifo_rf_din [DP-1:0];
    wire [DW-1:0] fifo_rf_r [DP-1:0];
    wire [DP-1:0] fifo_rf_en;
    wire wen = i_vld & i_rdy & i_clk_en;
    wire ren = o_vld & o_rdy & o_clk_en;
    wire [DP-1:0] rptr_vec_din; 
    wire [DP-1:0] rptr_vec_nxt;
    wire [DP-1:0] rptr_vec_r;
    wire [DP-1:0] wptr_vec_nxt;
    wire [DP-1:0] wptr_vec_r;
      if (DP == 1) begin:gen_wrptr_dp_1
          assign rptr_vec_nxt = 1'b1;
          assign wptr_vec_nxt = 1'b1;
      end
      else begin:gen_wrptr_dp_not_1
          assign rptr_vec_nxt =
            rptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                            (rptr_vec_r << 1);
          assign wptr_vec_nxt =
            wptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                            (wptr_vec_r << 1);
      end
e603_subsys_gnrl_dfflrs #(1)    rptr_vec_0_dfflrs  (ren, rptr_vec_nxt[0]     , rptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflrs #(1)    wptr_vec_0_dfflrs  (wen, wptr_vec_nxt[0]     , wptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
      if(DP>1) begin:gen_dp_gt1
e603_subsys_gnrl_dfflr  #(DP-1) rptr_vec_31_dfflr  (ren, rptr_vec_nxt[DP-1:1], rptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP-1) wptr_vec_31_dfflr  (wen, wptr_vec_nxt[DP-1:1], wptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
      end
    assign rptr_vec_din = ren ? rptr_vec_nxt : rptr_vec_r;
    wire [DP:0] i_vec;
    wire [DP:0] o_vec;
    wire [DP:0] vec_nxt;
    wire [DP:0] vec_r;
    wire vec_en = (ren ^ wen );
    assign vec_nxt = wen ? {vec_r[DP-1:0], 1'b1} : (vec_r >> 1);
e603_subsys_gnrl_dfflrs #(1)  vec_0_dfflrs     (vec_en, vec_nxt[0]     , vec_r[0]     ,     clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP) vec_31_dfflr     (vec_en, vec_nxt[DP:1], vec_r[DP:1],     clk, rst_n);// VPP_NO_REG_PARSE
    assign i_vec = {1'b0,vec_r[DP:1]};
    assign o_vec = {1'b0,vec_r[DP:1]};
  wire fifo_i_active;
  if (I_SUPPORT_RATIO == 0) begin : gen_i_no_ratio
    assign i_rdy = (~i_vec[DP-1]);
    assign fifo_i_active = 1'b0;
  end
  else begin: gen_i_ratio
    wire i_rdy_r_ena;
    wire i_rdy_r_nxt;
    wire i_rdy_r;
    wire i_need_updat;
    wire i_need_updat_r_set;
    wire i_need_updat_r_clr;
    wire i_need_updat_r_ena;
    wire i_need_updat_r_nxt;
    wire i_need_updat_r;
    assign i_need_updat = vec_en;
    assign i_need_updat_r_set = (i_need_updat && !i_clk_en);
    assign i_need_updat_r_clr = (i_need_updat_r && i_clk_en);
    assign i_need_updat_r_ena = i_need_updat_r_set || i_need_updat_r_clr;
    assign i_need_updat_r_nxt = i_need_updat_r_set;
e603_subsys_gnrl_dfflr  #(1) i_need_updat_r_dfflr    (i_need_updat_r_ena, i_need_updat_r_nxt, i_need_updat_r,     clk, rst_n);// VPP_NO_REG_PARSE
    assign i_rdy_r_ena = i_clk_en && (i_need_updat || i_need_updat_r);
    assign i_rdy_r_nxt = (vec_en) ? (~vec_nxt[DP]) : (~i_vec[DP-1]);
e603_subsys_gnrl_dfflrs  #(1) i_rdy_r_dfflrs    (i_rdy_r_ena, i_rdy_r_nxt, i_rdy_r,     clk, rst_n);// VPP_NO_REG_PARSE
    assign i_rdy = i_rdy_r;
    assign fifo_i_active = i_need_updat_r;
  end
    for (i=0; i<DP; i=i+1) begin:gen_fifo_rf
      assign fifo_rf_en[i] = wen & wptr_vec_r[i];
      if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_dffl   #(DW) fifo_rf_dffl  (fifo_rf_en[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      end
      else begin: rst_gen
e603_subsys_gnrl_dfflr  #(DW) fifo_rf_dfflr (fifo_rf_en[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      end
      assign fifo_rf_din[i] = fifo_rf_en[i] ? i_dat : fifo_rf_r[i];
    end
    integer j;
    wire [DW-1:0] mux_rdat;
    if(REG_OUT == 0) begin:gen_rdat_output
    reg [DW-1:0] mux_rdat_t;
        always @*
        begin : rd_port_PROC
          mux_rdat_t = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_t = mux_rdat_t | ({DW{rptr_vec_r[j]}} & fifo_rf_r[j]);
          end
        end
    assign mux_rdat = mux_rdat_t;
    if (O_SUPPORT_RATIO == 0) begin : gen_o_no_ratio
        assign o_dat = mux_rdat;
    end
    else begin: gen_o_ratio
        assign o_dat = mux_rdat & {DW{o_vld}};
    end
    end
    else begin:gen_rdat_flp_output
        reg [DW-1:0] mux_rdat_din;
        always @*
        begin : rd_port_PROC
          mux_rdat_din = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_din = mux_rdat_din | ({DW{rptr_vec_din[j]}} & fifo_rf_din[j]);
          end
        end
        wire mux_rdat_ena = 
                     (~o_vld) ? wen :
                     (vec_nxt[0] & ren);
e603_subsys_gnrl_dfflr #(DW) mux_rdat_dfflr  (mux_rdat_ena, mux_rdat_din, mux_rdat, clk, rst_n);// VPP_NO_REG_PARSE
    assign o_dat = mux_rdat;
    end
  wire fifo_o_active;
  if (O_SUPPORT_RATIO == 0) begin : gen_o_no_ratio
    assign o_vld = (o_vec[0]);
    assign fifo_o_active = 1'b0;
  end
  else begin : gen_o_ratio
    wire o_vld_r_ena;
    wire o_vld_r_nxt;
    wire o_vld_r;
    wire o_need_updat;
    wire o_need_updat_r_set;
    wire o_need_updat_r_clr;
    wire o_need_updat_r_ena;
    wire o_need_updat_r_nxt;
    wire o_need_updat_r;
    assign o_need_updat = vec_en;
    assign o_need_updat_r_set = (o_need_updat   && !o_clk_en);
    assign o_need_updat_r_clr = (o_need_updat_r &&  o_clk_en);
    assign o_need_updat_r_ena = o_need_updat_r_set || o_need_updat_r_clr;
    assign o_need_updat_r_nxt = o_need_updat_r_set;
e603_subsys_gnrl_dfflr  #(1) o_need_updat_r_dfflr    (o_need_updat_r_ena, o_need_updat_r_nxt, o_need_updat_r,     clk, rst_n);// VPP_NO_REG_PARSE
    assign o_vld_r_ena = o_clk_en && (o_need_updat || o_need_updat_r);
    assign o_vld_r_nxt = (vec_en) ? (vec_nxt[1]) : (o_vec[0]);
e603_subsys_gnrl_dfflr  #(1) o_vld_r_dfflr    (o_vld_r_ena, o_vld_r_nxt, o_vld_r,     clk, rst_n);// VPP_NO_REG_PARSE
    assign o_vld = o_vld_r;
    assign fifo_o_active = o_need_updat_r;
  end
  assign o_fifo_active =  i_vld || fifo_i_active || o_vld || fifo_o_active;
  end
endgenerate
endmodule
module e603_subsys_gnrl_loop_stck # (
  parameter PAYLOAD_NORST = 0,
    parameter DP = 4,
    parameter DW = 32
)(
    input  i_wen,
    input  o_ren,
    input  [DW-1:0] i_dat,
    output [DW-1:0] o_dat,
    input  clk,
    input  rst_n
);
  wire [DW-1:0] stck_rf_r [DP-1:0];
  wire [DP-1:0] stck_rf_en;
  wire [DP-1:0] i_vec;
  wire [DP-1:0] o_vec;
  wire [DP-1:0] vec_nxt;
  wire [DP-1:0] vec_r;
  wire vec_en = (o_ren ^ i_wen);
  assign vec_nxt =     o_ren ?
                   (vec_r[0] ? {1'b1,{DP-1{1'b0}}} : (vec_r >> 1)) :
                (vec_r[DP-1] ? {{DP-1{1'b0}},1'b1} : (vec_r << 1))
                             ;
e603_subsys_gnrl_dfflrs #(1)    vec_0_dfflrs(vec_en, vec_nxt[0]     , vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP-1) vec_dp_dfflr(vec_en, vec_nxt[DP-1:1], vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
  assign i_vec = vec_r; 
  assign o_vec = (vec_r == {{DP-1{1'b0}},1'b1}) ? {1'b1, {DP-1{1'b0}}}
                                                : (vec_r >> 1); 
  genvar i;
  generate 
    for (i=0; i<DP; i=i+1) begin:gen_stck_rf
      assign stck_rf_en[i] = i_wen & i_vec[i];      
      if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_dffl   #(DW) stck_rf_dffl  (stck_rf_en[i], i_dat, stck_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      end
      else begin: rst_gen
e603_subsys_gnrl_dfflr  #(DW) stck_rf_dfflr (stck_rf_en[i], i_dat, stck_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
      end
    end
  endgenerate
  integer j;
  reg [DW-1:0] mux_rdat;
  always @*
  begin : rd_port_PROC
    mux_rdat = {DW{1'b0}};
    for(j=0; j<DP; j=j+1) begin
      mux_rdat = mux_rdat | ({DW{o_vec[j]}} & stck_rf_r[j]);
    end
  end
  assign o_dat = mux_rdat;
endmodule
module e603_subsys_gnrl_cdc_buf
# (
  parameter PAYLOAD_NORST = 0,
  parameter I_ACTIVE_CUT_IVLD = 0,
  parameter DW = 32,
  parameter SYNC_DP = 2
) (
  input  i_clk,
  input  i_rst_n,
  input  i_vld,
  output i_rdy,
  input  [DW-1:0] i_dat,
  output i_cdc_buf_active,
  output o_cdc_buf_active,
  input  o_clk,
  input  o_rst_n,
  output o_vld,
  input  o_rdy,
  output [DW-1:0] o_dat
);
  wire tx_vld;
  wire tx_rdy;
  wire [DW-1:0] tx_dat;
  e603_subsys_gnrl_cdc_tx # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DW(DW),
    .SYNC_DP(SYNC_DP)
  ) u_cmd_cdc_tx(
    .i_vld  (i_vld),
    .i_rdy  (i_rdy),
    .i_dat  (i_dat),
    .o_vld  (tx_vld ),
    .o_rdy_a(tx_rdy ),
    .o_dat  (tx_dat),
    .clk    (i_clk),
    .rst_n  (i_rst_n)
  );
  e603_subsys_gnrl_cdc_rx # (
    .PAYLOAD_NORST(PAYLOAD_NORST),
    .DW(DW),
    .SYNC_DP(SYNC_DP)
   ) u_cmd_cdc_rx(
    .i_vld_a (tx_vld ),
    .i_rdy   (tx_rdy ),
    .i_dat   (tx_dat),
    .o_vld   (o_vld),
    .o_rdy   (o_rdy),
    .o_dat   (o_dat ),
    .clk    (o_clk),
    .rst_n  (o_rst_n)
  );
    generate 
        if(I_ACTIVE_CUT_IVLD == 1) begin: cut_ivld_gen
  assign i_cdc_buf_active = tx_vld;
        end
        else begin: no_cut_ivld_gen
  assign i_cdc_buf_active = i_vld  | tx_vld;
        end
    endgenerate
  assign o_cdc_buf_active = tx_rdy | o_vld;
endmodule
module e603_subsys_gnrl_2w1r_fifo # (
  parameter PAYLOAD_NORST = 0,
  parameter CUT_READY = 0,
  parameter MSKO = 0,
  parameter FIFO_REG_OUT = 0,
  parameter DP   = 8,
  parameter DW   = 32
) (
  input           i_vld0,
  input           i_vld1,
  output          i_rdy,
  input  [DW-1:0] i_dat0,
  input  [DW-1:0] i_dat1,
  output          o_vld,
  input           o_rdy,
  output [DW-1:0] o_dat,
  input           clk,
  input           rst_n
);
    wire [DW-1:0] fifo_rf_din [DP-1:0];
    wire [DW-1:0] fifo_rf_wdat [DP-1:0];
    wire [DW-1:0] fifo_rf_r [DP-1:0];
    wire [DP-1:0] fifo_rf_en0;
    wire [DP-1:0] fifo_rf_en1;
    wire [DP-1:0] fifo_rf_en;
    wire wen0 = i_vld0 & i_rdy;
    wire wen1 = i_vld1 & i_rdy;
    wire wen = (i_vld0 | i_vld1) & i_rdy;
    wire ren = o_vld & o_rdy;
    wire dual_wen = wen0 & wen1;
    wire [DP-1:0] rptr_vec_nxt;
    wire [DP-1:0] rptr_vec_din;
    wire [DP-1:0] rptr_vec_r;
    wire [DP-1:0] wptr_vec_nxt;
    wire [DP-1:0] wptr_vec_r;
    wire [DP-1:0] wptr_vec_r_lshift_1 = wptr_vec_r << 1;
    wire [DP-1:0] wptr0_vec_r = wptr_vec_r;
    wire [DP-1:0] wptr1_vec_r = wptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} : wptr_vec_r_lshift_1;
    assign rptr_vec_nxt =
          rptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                          (rptr_vec_r << 1);
    assign wptr_vec_nxt =
          wptr_vec_r[DP-1] ? (dual_wen ? {{DP-2{1'b0}}, 2'b10} : {{DP-1{1'b0}}, 1'b1}):
          wptr_vec_r[DP-2] ? (dual_wen ? {{DP-1{1'b0}}, 1'b1}  : wptr_vec_r_lshift_1):
                             (dual_wen ? (wptr_vec_r << 2)    : wptr_vec_r_lshift_1);
e603_subsys_gnrl_dfflrs #(1)    rptr_vec_0_dfflrs (ren, rptr_vec_nxt[0]     , rptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflrs #(1)    wptr_vec_0_dfflrs (wen, wptr_vec_nxt[0]     , wptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP-1) rptr_vec_31_dfflr (ren, rptr_vec_nxt[DP-1:1], rptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP-1) wptr_vec_31_dfflr (wen, wptr_vec_nxt[DP-1:1], wptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
    assign rptr_vec_din = ren  ? rptr_vec_nxt : rptr_vec_r;
    wire [DP:0] i_vec;
    wire [DP:0] o_vec;
    wire [DP:0] vec_nxt;
    wire [DP:0] vec_r;
    wire vec_en =
                 (~(   (~(ren | wen0 | wen1)) 
                      | (ren & (wen0 ^ wen1))  
                    ))
                ;
    assign vec_nxt =
                        ((~ren) & wen0 & wen1)  ? {vec_r[DP-2:0], 2'b11} :
                      (ren & (~wen0) & (~wen1)) ? (vec_r >> 1)
                                                : {vec_r[DP-1:0], 1'b1}
                                                ;
e603_subsys_gnrl_dfflrs #(1)  vec_0_dfflrs     (vec_en, vec_nxt[0]   , vec_r[0]   ,     clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP) vec_31_dfflr     (vec_en, vec_nxt[DP:1], vec_r[DP:1],     clk, rst_n);// VPP_NO_REG_PARSE
    assign i_vec = {1'b0,vec_r[DP:1]};
    assign o_vec = {1'b0,vec_r[DP:1]};
    genvar i;
    generate 
    assign i_rdy = (~i_vec[DP-2]) | ((~i_vec[DP-1]) & (~(i_vld0 & i_vld1)));
      for (i=0; i<DP; i=i+1) begin:gen_fifo_rf
        assign fifo_rf_en0[i] = ((wen0|wen1) & wptr0_vec_r[i]);
        assign fifo_rf_en1[i] = ((wen0&wen1) & wptr1_vec_r[i]);
        assign fifo_rf_en[i]  = fifo_rf_en0[i] | fifo_rf_en1[i];
        assign fifo_rf_wdat[i] = ({DW{fifo_rf_en0[i]}} & (wen0 ? i_dat0 : i_dat1))
                               | ({DW{fifo_rf_en1[i]}} & i_dat1)
                               ;
        if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_dffl   #(DW) fifo_rf_dffl  (fifo_rf_en[i],fifo_rf_wdat[i], fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
        end
        else begin: rst_gen
e603_subsys_gnrl_dfflr  #(DW) fifo_rf_dfflr (fifo_rf_en[i],fifo_rf_wdat[i], fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
        end
        assign fifo_rf_din[i] = fifo_rf_en[i] ? fifo_rf_wdat[i] : fifo_rf_r[i];
      end
    integer j;
    reg [DW-1:0] mux_rdat;
    if(FIFO_REG_OUT == 0) begin:gen_rdat_output
        always @*
        begin : rd_port_PROC
          mux_rdat = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat = mux_rdat | ({DW{rptr_vec_r[j]}} & fifo_rf_r[j]);
          end
        end
    end
    else begin:gen_rdat_flp_output
        reg [DW-1:0] mux_rdat_din;
        wire [DW-1:0] mux_rdat_r;
        always @*
        begin : rd_port_PROC
          mux_rdat_din = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_din = mux_rdat_din | ({DW{rptr_vec_din[j]}} & fifo_rf_din[j]);
          end
        end
e603_subsys_gnrl_dffr #(DW) mux_rdat_dffr  (mux_rdat_din, mux_rdat_r, clk, rst_n);// VPP_NO_REG_PARSE
        always @*
        begin : direct_assign
            mux_rdat = mux_rdat_r;
        end
    end
    endgenerate
    assign o_dat = mux_rdat;
    assign o_vld = (o_vec[0]);
endmodule
module e603_subsys_gnrl_cdc_pulse
# (
  parameter I_ACTIVE_CUT_IVLD = 0,
  parameter SYNC_DP = 2
) (
  input  i_clk,
  input  i_rst_n,
  input  i_pulse,
  output i_active,
  output o_active,
  input  o_clk,
  input  o_rst_n,
  output o_pulse
);
e603_subsys_gnrl_cdc_buf
# (
    .DW         (1      ),
    .I_ACTIVE_CUT_IVLD (I_ACTIVE_CUT_IVLD),
    .SYNC_DP    (SYNC_DP)
) u_gnrl_cdc_buf (
    .i_clk           (i_clk       ),
    .i_rst_n         (i_rst_n     ),
    .i_vld           (i_pulse     ),
    .i_rdy           (            ),
    .i_dat           (1'b0        ),
    .i_cdc_buf_active(i_active    ),
    .o_cdc_buf_active(o_active    ),
    .o_clk           (o_clk       ),
    .o_rst_n         (o_rst_n     ),
    .o_vld           (o_pulse     ),
    .o_rdy           (1'b1        ),
    .o_dat           (            )
);
endmodule
module e603_subsys_gnrl_cdc_fifo #(
  parameter PAYLOAD_NORST = 0,
  parameter SMALL_DP_EN    = 0,
  parameter SMALL_DP       = 6,
  parameter SMALL_DP_PTR_W = 3,
  parameter DP   = 5,
  parameter DP_PTR_W   = 3,
  parameter DW   = 32,
  parameter SYNC_DP = 2
) (
  input  i_clk,
  input  i_rst_n,
  input  i_vld,
  output i_rdy,
  input  [DW-1:0] i_dat,
  output i_cdc_fifo_active,
  output o_cdc_fifo_active,
  input  o_clk,
  input  o_rst_n,
  output o_vld,
  input  o_rdy,
  output [DW-1:0] o_dat
);
  wire          wr   ;
  wire [DW-1:0] wdata;
  wire          full ;
  wire          rd   ;
  wire [DW-1:0] rdata;
  wire          empty;
  wire          w_empty;
  e603_subsys_gnrl_async_fifo #(.DW(DW), .DP(DP),  .DP_PTR_W(DP_PTR_W), .SYNC_DP(SYNC_DP), 
                               .SMALL_DP_EN(SMALL_DP_EN),
       .PAYLOAD_NORST(PAYLOAD_NORST),
                               .SMALL_DP(SMALL_DP),  .SMALL_DP_PTR_W(SMALL_DP_PTR_W))
  u_a_fifo (
    .wclk     (i_clk),
    .wrst_n   (i_rst_n),
    .wr       (wr),
    .wdata    (wdata),
    .wwmk     (),
    .full     (full),
    .w_empty  (w_empty),
    .rclk     (o_clk),
    .rrst_n   (o_rst_n),
    .rd       (rd),
    .rdata    (rdata),
    .rwmk     (),
    .empty    (empty)
  );
  assign i_rdy = ~full;
  assign wr = i_vld & i_rdy;
  assign wdata = i_dat;
  assign o_vld = ~empty;
  assign rd = o_vld & o_rdy;
  assign o_dat = rdata;
  assign i_cdc_fifo_active = (~w_empty);
  assign o_cdc_fifo_active = ~empty;
endmodule
module e603_subsys_gnrl_data_mux # (
  parameter DW = 8,
  parameter N  = 2,
  parameter SW = N<=1 ? 1 : N<=2**0 ? 0 : N<=2**1 ? 1 : N<=2**2 ? 2 : N<=2**3 ? 3 : N<=2**4 ? 4 : N<=2**5 ? 5 : N<=2**6 ? 6 : N<=2**7 ? 7 : N<=2**8 ? 8 : N<=2**9 ? 9 : N<=2**10 ? 10 : N<=2**11 ? 11 : N<=2**12 ? 12 : N<=2**13 ? 13 : N<=2**14 ? 14 : N<=2**15 ? 15 : N<=2**16 ? 16 : N<=2**17 ? 17 : N<=2**18 ? 18 : N<=2**19 ? 19 : N<=2**20 ? 20 : N<=2**21 ? 21 : N<=2**22 ? 22 : N<=2**23 ? 23 : N<=2**24 ? 24 : N<=2**25 ? 25 : N<=2**26 ? 26 : N<=2**27 ? 27 : N<=2**28 ? 28 : N<=2**29 ? 29 : N<=2**30 ? 30 : N<=2**31 ? 31 : 32
)(
  output   [DW-1:0] out_data,
  input  [N*DW-1:0] in_data,
  input    [SW-1:0] sel
);
  wire [DW-1:0] in_data_xy [N-1:0];
  wire  [N-1:0] in_data_yx [DW-1:0];
  wire  [N-1:0] in_data_mask;
  genvar gvi, gvj;
  generate
  for (gvi=0; gvi<N; gvi=gvi+1) begin: GEN_in_data_xy
    assign in_data_xy[gvi] = in_data[gvi*DW +: DW];
    assign in_data_mask[gvi] = (gvi[SW-1:0] == sel);
    for (gvj=0; gvj<DW; gvj=gvj+1) begin: GEN_in_data_yx
      assign in_data_yx[gvj][gvi] = in_data_xy[gvi][gvj];
    end 
  end 
  for (gvi=0; gvi<DW; gvi=gvi+1) begin: GEN_out_data
    assign out_data[gvi] = |(in_data_mask & in_data_yx[gvi]);
  end 
  endgenerate
endmodule
module e603_subsys_gnrl_mem_line #(
  parameter DW = 8
)(
  input           clk,
  input           rst_n,
  input           wr,
  input  [DW-1:0] wdata,
  output [DW-1:0] mem
);
e603_subsys_gnrl_dfflr #(DW) mem_dfflr (wr, wdata, mem, clk, rst_n);// VPP_NO_REG_PARSE
endmodule
module e603_subsys_gnrl_async_mem_line #(
  parameter PAYLOAD_NORST = 0,
  parameter DW = 8
)(
  input           clk,
  input           rst_n,
  input           wr,
  input  [DW-1:0] wdata,
  output [DW-1:0] mem
);
      generate
        if(PAYLOAD_NORST == 1) begin: payload_norst
      e603_subsys_gnrl_cdc_dffl  #(DW) mem_dffl  (wr, wdata, mem, clk, rst_n);  // VPP_NO_REG_PARSE
        end
        else begin: payload_rst
      e603_subsys_gnrl_cdc_dfflr #(DW) mem_dfflr (wr, wdata, mem, clk, rst_n);  // VPP_NO_REG_PARSE
        end
      endgenerate
endmodule
module e603_subsys_gnrl_hsk_arbt # (
  parameter DW = 64,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_NUM = 4,
  parameter ARBT_PTR_W = 2
) (
  output          arbt_active,
  input           clk_en,
  output          o_valid,
  input           o_ready,
  output [DW-1:0] o_data,
  output          o_first,
  output          o_last,
  output [ARBT_NUM*1-1:0]     i_bus_ready,
  input  [ARBT_NUM*1-1:0]     i_bus_valid,
  input  [ARBT_NUM*DW-1:0]    i_bus_data,
  input  [ARBT_NUM-1:0]       i_bus_first,
  input  [ARBT_NUM-1:0]       i_bus_last,
  input  [ARBT_NUM*1-1:0]     i_bus_sel_vec,
  output [ARBT_NUM*1-1:0]     o_bus_sel_vec,
  input  clk,
  input  rst_n
  );
  localparam ARBT_SCHEME_PRIORITY  = 0;
  localparam ARBT_SCHEME_RROBIN    = 1;
  localparam ARBT_SCHEME_DIRECT_SEL_1HOT = 2;
  localparam ARBT_SCHEME_DIRECT_SEL_PRIORITY = 3;
  localparam ARBT_SCHEME_RROBIN4   = 4;
  wire rrobin_active;
  wire [ARBT_NUM-1:0] burst_mask_r;
  wire [ARBT_NUM*1-1:0] i_bus_sel_vec_pos;
  wire [ARBT_NUM*1-1:0] i_bus_ready_pos;
  wire [ARBT_NUM*1-1:0] i_bus_valid_pos;
genvar i;
generate 
  if(ARBT_NUM == 1) begin:gen_arbt_num_eq_1
    assign i_bus_ready   = o_ready    ;
    assign o_valid       = i_bus_valid;
    assign o_data        = i_bus_data;
    assign o_first       = i_bus_first;
    assign o_last        = i_bus_last;
    assign rrobin_active = 1'b0;
    assign burst_mask_r = {ARBT_NUM{1'b0}};
    assign o_bus_sel_vec = 1'b1;
  end
  else begin:gen_arbt_num_gt_1
    integer j;
    wire [ARBT_NUM-1:0] i_bus_grt_vec;
    wire [ARBT_NUM-1:0] i_bus_sel;
    wire [DW-1:0] i_data[ARBT_NUM-1:0];
    wire [1-1:0]  i_first[ARBT_NUM-1:0];
    wire [1-1:0]  i_last [ARBT_NUM-1:0];
    reg [DW-1:0] sel_o_data;
    reg          sel_o_first;
    reg          sel_o_last;
    assign o_bus_sel_vec = i_bus_sel;
    wire arbt_ena;
    wire [ARBT_NUM-1:0] burst_mask_nxt;
    wire burst_mask_ena;
    wire burst_mask_set;
    wire burst_mask_clr;
    assign burst_mask_set = o_first & arbt_ena;
    assign burst_mask_clr = (|burst_mask_r) & o_last & arbt_ena;
    assign burst_mask_ena = clk_en & (burst_mask_set | burst_mask_clr);
    assign burst_mask_nxt = burst_mask_clr ? {ARBT_NUM{1'b0}} : (~i_bus_sel); 
e603_subsys_gnrl_dfflr #(ARBT_NUM) burst_mask_dfflr (burst_mask_ena, burst_mask_nxt, burst_mask_r, clk, rst_n);// VPP_NO_REG_PARSE
    assign i_bus_valid_pos   = (~burst_mask_r) & i_bus_valid;
    assign i_bus_ready       = (~burst_mask_r) & i_bus_ready_pos;
    assign i_bus_sel_vec_pos = (~burst_mask_r) & i_bus_sel_vec;
    for(i = 0; i < ARBT_NUM; i = i+1)
    begin:gen_distract
      assign i_data [i] = i_bus_data[(i+1)*DW-1 : i*DW    ];
      assign i_first[i] = i_bus_first[(i+1)*1-1 : i*1    ];
      assign i_last [i] = i_bus_last [(i+1)*1-1 : i*1    ];
      assign i_bus_ready_pos[i] = i_bus_grt_vec[i] & o_ready;
    end
    assign arbt_ena = o_valid & o_ready;
    if(ARBT_SCHEME == ARBT_SCHEME_PRIORITY) begin:gen_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_grt_vec[i] =  1'b1;
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_valid_pos[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_grt_vec[i] =  ~(|i_bus_valid_pos[i-1:0]);
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_valid_pos[i];
        end
      end
      assign o_valid = |i_bus_valid_pos;
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN) begin:gen_rrobin_arbt
     e603_subsys_gnrl_rrobin # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin(
       .rrobin_active (rrobin_active),
       .grt_vec  (i_bus_grt_vec),
       .req_vec  (i_bus_valid_pos),
       .arbt_ena (arbt_ena & clk_en),
       .clk      (clk),
       .rst_n    (rst_n)
     );
     assign i_bus_sel = i_bus_grt_vec;
     assign o_valid = |i_bus_valid_pos;
   end
   else begin: gen_no_rrobin
     assign rrobin_active = 1'b0;
   end
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_1HOT) begin:gen_indic_arbt
     assign i_bus_grt_vec = i_bus_sel_vec_pos;
     assign i_bus_sel = i_bus_grt_vec;
     assign o_valid = |(i_bus_valid_pos & i_bus_sel_vec_pos);
   end
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_PRIORITY) begin:gen_indic_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_grt_vec[i] =  1'b1;
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_sel_vec_pos[i];
        end
        else if(i==(ARBT_NUM-1)) begin: gen_i_is_n
          assign i_bus_grt_vec[i] =  ~(|i_bus_sel_vec_pos[i-1:0]);
          assign i_bus_sel[i] = i_bus_grt_vec[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_grt_vec[i] =  ~(|i_bus_sel_vec_pos[i-1:0]);
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_sel_vec_pos[i];
        end
      end
      assign o_valid = |(i_bus_valid_pos & i_bus_sel);
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN4) begin:gen_rbin4_arbt
      e603_subsys_gnrl_rbin4 # (
          .ARBT_NUM(ARBT_NUM)
      )u_e603_subsys_gnrl_rbin4(
        .grt_vec  (i_bus_grt_vec),
        .req_vec  (i_bus_sel_vec_pos),
        .arbt_ena (arbt_ena & clk_en & (~burst_mask_set)),
        .rbin4_active (),
        .clk      (clk),
        .rst_n    (rst_n)
      );
      assign i_bus_sel = i_bus_grt_vec & i_bus_sel_vec_pos;
      assign o_valid = |(i_bus_valid_pos & i_bus_sel);
   end
    always @ (*) begin : sel_o_ready_PROC
      sel_o_data  = {DW  {1'b0}};
      sel_o_first = 1'b0;
      sel_o_last  = 1'b0;
      for(j = 0; j < ARBT_NUM; j = j+1) begin
        sel_o_data  = sel_o_data  | ({DW{i_bus_sel[j]}} & i_data [j]);
        sel_o_first = sel_o_first | (    i_bus_sel[j]   & i_first[j]);
        sel_o_last  = sel_o_last  | (    i_bus_sel[j]   & i_last [j]);
      end
    end
    assign o_data  = sel_o_data;
    assign o_first = sel_o_first;
    assign o_last  = sel_o_last;
  end
  endgenerate 
  assign arbt_active = (|i_bus_valid) | rrobin_active;
endmodule
module e603_subsys_gnrl_hsk_arbt_1cycle # (
  parameter DW = 64,
  parameter ARBT_SCHEME = 3,
  parameter ARBT_NUM = 4,
  parameter ARBT_PTR_W = 2
) (
  output          arbt_active,
  input           clk_en,
  output          o_valid,
  input           o_ready,
  output [DW-1:0] o_data,
  output [ARBT_NUM*1-1:0]     i_bus_ready,
  input  [ARBT_NUM*1-1:0]     i_bus_valid,
  input  [ARBT_NUM*1-1:0]     i_bus_busy,
  input  [ARBT_NUM*DW-1:0]    i_bus_data,
  input                       i_bus_grt_rply,
  input  [ARBT_NUM*1-1:0]     i_bus_sel_vec,
  output [ARBT_NUM*1-1:0]     o_bus_sel_vec,
  input  clk,
  input  rst_n
  );
  localparam ARBT_SCHEME_PRIORITY  = 0;
  localparam ARBT_SCHEME_RROBIN    = 1;
  localparam ARBT_SCHEME_DIRECT_SEL_1HOT = 2;
  localparam ARBT_SCHEME_DIRECT_SEL_PRIORITY = 3;
  localparam ARBT_SCHEME_RROBIN4   = 4;
  localparam ARBT_SCHEME_RROBIN_DA = 6;
  wire rrobin_active;
  wire [ARBT_NUM*1-1:0] i_bus_sel_vec_pos;
  wire [ARBT_NUM*1-1:0] i_bus_ready_pos;
  wire [ARBT_NUM*1-1:0] i_bus_valid_pos;
genvar i;
generate 
  if(ARBT_NUM == 1) begin:gen_arbt_num_eq_1
    assign i_bus_ready   = o_ready    ;
    assign o_valid       = i_bus_valid;
    assign o_data        = i_bus_data;
    assign rrobin_active = 1'b0;
    assign o_bus_sel_vec = 1'b1;
  end
  else begin:gen_arbt_num_gt_1
    integer j;
    wire [ARBT_NUM-1:0] i_bus_grt_vec;
    wire [ARBT_NUM-1:0] i_bus_sel;
    wire [DW-1:0] i_data[ARBT_NUM-1:0];
    reg [DW-1:0] sel_o_data;
    assign o_bus_sel_vec = i_bus_sel;
    wire arbt_ena;
    assign i_bus_valid_pos   = i_bus_valid;
    assign i_bus_ready       = i_bus_ready_pos;
    assign i_bus_sel_vec_pos = i_bus_sel_vec;
    for(i = 0; i < ARBT_NUM; i = i+1)
    begin:gen_distract
      assign i_data [i] = i_bus_data[(i+1)*DW-1 : i*DW    ];
      assign i_bus_ready_pos[i] = i_bus_grt_vec[i] & o_ready;
    end
    assign arbt_ena = o_valid & o_ready;
    if(ARBT_SCHEME == ARBT_SCHEME_PRIORITY) begin:gen_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_grt_vec[i] =  1'b1;
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_valid_pos[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_grt_vec[i] =  ~(|i_bus_valid_pos[i-1:0]);
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_valid_pos[i];
        end
      end
      assign o_valid = |i_bus_valid_pos;
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN) begin:gen_rrobin_arbt
    wire rrobin_arbt_ena = clk_en & o_ready;
     e603_subsys_gnrl_rrobin_1cycle # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin(
       .rrobin_active (rrobin_active),
       .grt_vec  (i_bus_grt_vec),
       .req_vec  (i_bus_valid_pos),
       .arbt_ena (rrobin_arbt_ena),
       .clk      (clk),
       .rst_n    (rst_n)
     );
     assign i_bus_sel = i_bus_grt_vec;
     assign o_valid = |i_bus_valid_pos;
   end
   else if(ARBT_SCHEME == ARBT_SCHEME_RROBIN_DA) begin:gen_rrobin_da_arbt
    wire rrobin_arbt_ena = clk_en & o_ready;
     e603_subsys_gnrl_rrobin_1cycle_da # (
         .ARBT_NUM(ARBT_NUM)
     )u_e603_subsys_gnrl_rrobin(
       .rrobin_active (rrobin_active),
       .grt_vec  (i_bus_grt_vec),
       .buz_vec  (i_bus_busy),
       .req_vec  (i_bus_valid_pos),
       .arbt_ena (rrobin_arbt_ena),
       .arbt_rply(i_bus_grt_rply),
       .clk      (clk),
       .rst_n    (rst_n)
     );
     assign i_bus_sel = i_bus_grt_vec;
     assign o_valid = |i_bus_valid_pos;
   end
   else begin: gen_no_rrobin
     assign rrobin_active = 1'b0;
   end
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_1HOT) begin:gen_indic_arbt
     assign i_bus_grt_vec = i_bus_sel_vec_pos;
     assign i_bus_sel = i_bus_grt_vec;
     assign o_valid = |(i_bus_valid_pos & i_bus_sel_vec_pos);
   end
   if(ARBT_SCHEME == ARBT_SCHEME_DIRECT_SEL_PRIORITY) begin:gen_indic_priorty_arbt
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:gen_priroty_grt_vec
        if(i==0) begin: gen_i_is_0
          assign i_bus_grt_vec[i] =  1'b1;
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_sel_vec_pos[i];
        end
        else if(i==(ARBT_NUM-1)) begin: gen_i_is_n
          assign i_bus_grt_vec[i] =  ~(|i_bus_sel_vec_pos[i-1:0]);
          assign i_bus_sel[i] = i_bus_grt_vec[i];
        end
        else begin:gen_i_is_not_0
          assign i_bus_grt_vec[i] =  ~(|i_bus_sel_vec_pos[i-1:0]);
          assign i_bus_sel[i] = i_bus_grt_vec[i] & i_bus_sel_vec_pos[i];
        end
      end
      assign o_valid = |(i_bus_valid_pos & i_bus_sel);
    end
   if(ARBT_SCHEME == ARBT_SCHEME_RROBIN4) begin:gen_rbin4_arbt
      e603_subsys_gnrl_rbin4 # (
          .ARBT_NUM(ARBT_NUM)
      )u_e603_subsys_gnrl_rbin4(
        .grt_vec  (i_bus_grt_vec),
        .req_vec  (i_bus_sel_vec_pos),
        .rbin4_active (),
        .arbt_ena (clk_en),
        .clk      (clk),
        .rst_n    (rst_n)
      );
      assign i_bus_sel = i_bus_grt_vec & i_bus_sel_vec_pos;
      assign o_valid = |(i_bus_valid_pos & i_bus_sel);
   end
    always @ (*) begin : sel_o_ready_PROC
      sel_o_data  = {DW  {1'b0}};
      for(j = 0; j < ARBT_NUM; j = j+1) begin
        sel_o_data  = sel_o_data  | ({DW{i_bus_sel[j]}} & i_data [j]);
      end
    end
    assign o_data  = sel_o_data;
  end
  endgenerate 
  assign arbt_active = (|i_bus_valid) | rrobin_active;
endmodule
module e603_subsys_gnrl_xshft_rng (clk, rst_n, load, seed, en, rnd);
  localparam DW = 32;
  localparam [DW-1:0] INIT = 32'h0000_1208;
  input           clk;
  input           rst_n;
  input           load;
  input  [DW-1:0] seed;
  input           en;
  output [DW-1:0] rnd;
  wire [DW-1:0] xs_1 = rnd ^ (rnd >> 13);
  wire [DW-1:0] xs_2 = xs_1 ^ (xs_1 << 3);
  wire [DW-1:0] xs_3 = xs_2 ^ (xs_2 >> 17);
  wire          rnd_ena;
  wire [DW-1:0] rnd_nxt;
  assign rnd_ena = load | en;
  assign rnd_nxt = load ? seed : xs_3;
e603_subsys_gnrl_dfflrs #(DW,INIT) rnd_dfflr(rnd_ena, rnd_nxt, rnd, clk, rst_n);// VPP_NO_REG_PARSE
endmodule 
`include "global.v"
module e603_subsys_gnrl_cdc_rx
# (
  parameter PAYLOAD_NORST = 0,
  parameter READY_THROUGH = 0,
  parameter DW = 32,
  parameter SYNC_DP = 2
) (
  input  i_vld_a, 
  output i_rdy, 
  input  [DW-1:0] i_dat,
  output o_vld, 
  input  o_rdy, 
  output [DW-1:0] o_dat,
  input  clk,
  input  rst_n 
);
wire i_vld_sync;
e603_subsys_gnrl_sync #(.DP(SYNC_DP), .DW(1)) u_i_vld_sync (
     .clk   (clk),
     .rst_n (rst_n),
     .din_a (i_vld_a),
     .dout  (i_vld_sync)
    );
wire i_vld_sync_r;
e603_subsys_gnrl_dffr #(1) i_vld_sync_dffr(i_vld_sync, i_vld_sync_r, clk, rst_n);// VPP_NO_REG_PARSE
wire i_vld_sync_nedge = (~i_vld_sync) & i_vld_sync_r;
wire buf_rdy;
wire i_rdy_r;
wire buf_dat_ena;
wire i_rdy_set;
generate
  if(READY_THROUGH == 0) begin: no_ready_through_gen
    assign i_rdy_set = buf_rdy & i_vld_sync 
                 & (~i_rdy_r)
                 ;
    assign buf_dat_ena = i_rdy_set;
  end
  else begin: ready_through_gen
    assign i_rdy_set = i_vld_sync 
               & o_vld & o_rdy
               ;
    assign buf_dat_ena = (~i_rdy_r) & buf_rdy & i_vld_sync;
  end
endgenerate
wire i_rdy_clr = i_vld_sync_nedge;
wire i_rdy_ena = i_rdy_set |   i_rdy_clr;
wire i_rdy_nxt = i_rdy_set | (~i_rdy_clr);
e603_subsys_gnrl_cdc_dfflr #(1) i_rdy_gnrl_cdc_dfflr(i_rdy_ena, i_rdy_nxt, i_rdy_r, clk, rst_n); // VPP_NO_REG_PARSE
assign i_rdy = i_rdy_r;
wire buf_vld_r;
wire [DW-1:0] buf_dat_r;
generate
    if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_cdc_dffl  #(DW) buf_dat_gnrl_cdc_dest_dffl (buf_dat_ena, i_dat, buf_dat_r, clk, rst_n); // VPP_NO_REG_PARSE
    end
    else begin: rst_gen
e603_subsys_gnrl_cdc_dfflr #(DW) buf_dat_gnrl_cdc_dest_dfflr(buf_dat_ena, i_dat, buf_dat_r, clk, rst_n); // VPP_NO_REG_PARSE
    end
endgenerate
wire buf_vld_set = buf_dat_ena;
wire buf_vld_clr = o_vld & o_rdy;
wire buf_vld_ena = buf_vld_set | buf_vld_clr;
wire buf_vld_nxt = buf_vld_set | (~buf_vld_clr);
e603_subsys_gnrl_dfflr #(1) buf_vld_dfflr(buf_vld_ena, buf_vld_nxt, buf_vld_r, clk, rst_n);// VPP_NO_REG_PARSE
assign buf_rdy = (~buf_vld_r);
assign o_vld = buf_vld_r;
assign o_dat = buf_dat_r;
endmodule 
module e603_subsys_gnrl_cdc_ack_channel
# (
  parameter SYNC_DP = 2
) (
  input  req_a, 
  output ack_o, 
  output req_o, 
  input  clk,
  input  rst_n 
);
  e603_subsys_gnrl_cdc_rx # (
     .READY_THROUGH(1),
     .DW      (1),
     .SYNC_DP (SYNC_DP)
   ) u_cdc_ack_channel (
  .i_vld_a (req_a), 
  .i_rdy   (ack_o), 
  .i_dat   (1'b0),
  .o_vld   (req_o), 
  .o_rdy   (1'b1), 
  .o_dat   (),
  .clk     (clk),
  .rst_n   (rst_n)
);
endmodule
`include "global.v"
module e603_subsys_gnrl_async_fifo_ctl # (
  parameter DP = 4,
  parameter DP_PTR_W = 2,
  parameter WWMK = 1,
  parameter RWMK = 1,
  parameter SYNC_DP = 2,
  parameter        AW = (DP <= 1) ? 1 : DP_PTR_W 
)(
  input           wclk,
  input           wrst_n,
  input           wr,
  output          wwmk,
  output          full,
  output          w_empty,
  output [AW-1:0] waddr,
  input           rclk,
  input           rrst_n,
  input           rd,
  output          rwmk,
  output          empty,
  output [AW-1:0] raddr,
  output          r_cs
);
  localparam [AW:0] PTR_START = {{1'b1},{(AW){1'b0}}} - DP;
  localparam [AW:0] PTR_END   = (~PTR_START);
  localparam [AW:0] PTR_START_G = bin2gray(PTR_START);
  wire   [AW:0] rptr_g_wclk;
  wire          safe_wr;
  wire   [AW:0] wptr_nxt, wptr_g_nxt;
  wire [AW-1:0] waddr_nxt;
  wire   [AW:0] wptr_din, wptr_g_din;
  wire [AW-1:0] waddr_din;
  wire   [AW:0] wptr;
  wire   [AW:0] wptr_g;
  wire   [AW:0] rptr_wclk;
  wire [AW-1:0] raddr_wclk;
  wire          wroll_over;
  wire   [AW:0] wwmk_lmt;
  wire   [AW:0] wptr_g_rclk;
  wire          safe_rd;
  wire   [AW:0] rptr_nxt, rptr_g_nxt;
  wire   [AW:0] rptr_din, rptr_g_din;
  wire [AW-1:0] raddr_din;
  wire   [AW:0] rptr;
  wire   [AW:0] rptr_g;
  wire   [AW:0] wptr_rclk;
  wire [AW-1:0] waddr_rclk;
  wire          rroll_over;
  wire   [AW:0] rwmk_lmt;
  e603_subsys_gnrl_sync #(
  .DW(AW+1),
  .RST_VAL(PTR_START_G),
  .DP(SYNC_DP))
  U_rptr_g_wclk_sync (
  .clk(wclk),
  .rst_n(wrst_n),
  .din_a(rptr_g),
  .dout(rptr_g_wclk)
  );
  e603_subsys_gnrl_sync #(
  .DW(AW+1),
  .RST_VAL(PTR_START_G),
  .DP(SYNC_DP))
  U_wptr_g_rclk_sync (
  .clk(rclk),
  .rst_n(rrst_n),
  .din_a(wptr_g),
  .dout(wptr_g_rclk)
  );
  assign safe_wr = wr & (~full);
  assign wptr_nxt   = ((wptr == PTR_END) ? PTR_START : wptr + ({(AW+1){1'b1}} >> (AW+1-1)));
  assign wptr_g_nxt = bin2gray(wptr_nxt);
  assign waddr_nxt  = ptr2addr(wptr_nxt);
  assign wptr_din   = safe_wr ? wptr_nxt : wptr;
  assign wptr_g_din = bin2gray(wptr_din);
  assign waddr_din  = ptr2addr(wptr_din);
  assign wptr = gray2bin(wptr_g);
e603_subsys_gnrl_dfflrs #(AW+1, PTR_START_G) wptr_g_dfflrs (safe_wr, wptr_g_nxt, wptr_g, wclk, wrst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(AW)                waddr_dfflr   (safe_wr, waddr_nxt, waddr, wclk, wrst_n);// VPP_NO_REG_PARSE
  assign rptr_wclk = gray2bin(rptr_g_wclk);
  assign raddr_wclk = ptr2addr(rptr_wclk);
  assign wroll_over = (wptr_g_din[AW] ^ rptr_g_wclk[AW]);
  wire full_nxt;
  assign full_nxt = wroll_over & (waddr_din == raddr_wclk);
e603_subsys_gnrl_dffr #(1) full_dffr (full_nxt, full, wclk, wrst_n);// VPP_NO_REG_PARSE
  wire w_empty_nxt;
  assign w_empty_nxt = (~wroll_over) & (waddr_din == raddr_wclk);
e603_subsys_gnrl_dffrs #(1, 1'b1) w_empty_dffrs (w_empty_nxt, w_empty, wclk, wrst_n);// VPP_NO_REG_PARSE
  assign wwmk_lmt = wroll_over ? {1'b0, raddr_wclk} - (DP[AW:0]-WWMK[AW:0])
                               : {1'b0, raddr_wclk} + WWMK[AW:0];
  wire wwmk_nxt;
  assign wwmk_nxt = ({1'b0, waddr_din} >= wwmk_lmt) | (wroll_over & wwmk_lmt[AW]);
e603_subsys_gnrl_dffr #(1) wwmk_dffr (wwmk_nxt, wwmk, wclk, wrst_n);// VPP_NO_REG_PARSE
  assign safe_rd = rd & (~empty);
  wire empty_din;
  assign r_cs = (~empty_din) & (empty | rd);
  assign rptr_nxt   = ((rptr == PTR_END) ? PTR_START : rptr + ({(AW+1){1'b1}} >> (AW+1-1)));
  assign rptr_g_nxt = bin2gray(rptr_nxt);
  assign rptr_din   = safe_rd ? rptr_nxt : rptr;
  assign rptr_g_din = bin2gray(rptr_din);
  assign raddr_din  = ptr2addr(rptr_din);
  assign rptr = gray2bin(rptr_g);
e603_subsys_gnrl_dfflrs #(AW+1, PTR_START_G) rptr_g_dfflrs (safe_rd, rptr_g_nxt, rptr_g, rclk, rrst_n);// VPP_NO_REG_PARSE
  assign raddr = raddr_din;
  assign wptr_rclk = gray2bin(wptr_g_rclk);
  assign waddr_rclk = ptr2addr(wptr_rclk);
  assign rroll_over = (rptr_g_din[AW] ^ wptr_g_rclk[AW]);
  wire empty_nxt;
  assign empty_nxt = (~rroll_over) & (raddr_din == waddr_rclk);
e603_subsys_gnrl_dffrs #(1, 1'b1) empty_dffrs (empty_nxt, empty, rclk, rrst_n);// VPP_NO_REG_PARSE
  assign empty_din = empty_nxt;
  assign rwmk_lmt = rroll_over ? {1'b0, waddr_rclk} + (DP[AW:0]-RWMK[AW:0])
                               : {1'b0, waddr_rclk} - RWMK[AW:0];
  wire rwmk_nxt;
  assign rwmk_nxt = ({1'b0, raddr_din} <= rwmk_lmt) & (rroll_over | (~rwmk_lmt[AW]));
e603_subsys_gnrl_dffrs #(1, 1'b1) rwmk_dffrs (rwmk_nxt, rwmk, rclk, rrst_n);// VPP_NO_REG_PARSE
  function automatic [AW:0] bin2gray;
    input [AW:0] bin;
    bin2gray = bin ^ (bin>>1);
  endfunction
  function automatic [AW:0] gray2bin;
    input [AW:0] gray;
    integer i;
    for (i=0; i<AW+1; i=i+1) begin
      gray2bin[i] = (^(gray>>i));
    end
  endfunction
  function automatic [AW-1:0] ptr2addr;
    input [AW:0] ptr;
    ptr2addr = ptr[AW] ? ptr[AW-1:0] : (ptr[AW-1:0] - PTR_START[AW-1:0]);
  endfunction
endmodule 
module e603_subsys_gnrl_async_fifo #(
  parameter PAYLOAD_NORST    = 0,
  parameter SMALL_DP_EN    = 0,
  parameter SMALL_DP       = 6,
  parameter SMALL_DP_PTR_W = 3,
  parameter DW = 4,
  parameter DP = 4,
  parameter DP_PTR_W = 2,
  parameter WWMK = 1,
  parameter RWMK = 1,
  parameter SYNC_DP = 2 
)(
  input           wclk,
  input           wrst_n,
  input           wr,
  input  [DW-1:0] wdata,
  output          wwmk,
  output          full,
  output          w_empty,
  input           rclk,
  input           rrst_n,
  input           rd,
  output [DW-1:0] rdata,
  output          rwmk,
  output          empty
);
  localparam I_DP       = SMALL_DP_EN ? SMALL_DP       : (DP < 8 ) ? 8 : DP;
  localparam I_DP_PTR_W = SMALL_DP_EN ? SMALL_DP_PTR_W : (DP < 8 ) ? 3 : DP_PTR_W;
  localparam AW = I_DP_PTR_W;
  wire [AW-1:0] waddr, raddr;
 wire r_cs;
  e603_subsys_gnrl_async_fifo_ctl #(
  .DP(I_DP),
  .DP_PTR_W(I_DP_PTR_W),
  .WWMK(WWMK),
  .RWMK(RWMK),
  .SYNC_DP(SYNC_DP))
  U_ctl (
  .wclk(wclk),
  .wrst_n(wrst_n),
  .wr(wr),
  .full(full),
  .wwmk(wwmk),
  .waddr(waddr),
  .rclk(rclk),
  .rrst_n(rrst_n),
  .rd(rd),
  .empty(empty),
  .rwmk(rwmk),
  .raddr(raddr),
  .r_cs(r_cs),
  .w_empty(w_empty)
  );
  e603_subsys_gnrl_async_sdp_ram #(
  .PAYLOAD_NORST(PAYLOAD_NORST),
  .DW(DW),
  .DP(I_DP),
  .DP_PTR_W(AW),
  .REG_OUT(1))
  U_ram (
  .wclk(wclk),
  .wrst_n(wrst_n),
  .wr(wr),
  .waddr(waddr),
  .wdata(wdata),
  .rclk(rclk),
  .rrst_n(rrst_n),
  .rd(r_cs),
  .raddr(raddr),
  .rdata(rdata)
  );
endmodule 
`include "global.v"
module e603_subsys_gnrl_sdp_ram #(
  parameter DW = 8,
  parameter DP = 4,
  parameter DP_PTR_W = 2,
  parameter REG_OUT = 1,
  parameter AW = (DP <= 1) ? 1 : DP_PTR_W
)(
  input           wclk,
  input           wrst_n,
  input           wr,
  input  [AW-1:0] waddr,
  input  [DW-1:0] wdata,
  input           rclk,
  input           rrst_n,
  input           rd,
  input  [AW-1:0] raddr,
  output [DW-1:0] rdata
);
  wire    [DP-1:0] wword_line, rword_line;
  wire [DP*DW-1:0] mem;
  wire    [DW-1:0] rdata_int;
  genvar gvi;
  generate
  for (gvi=0; gvi<DP; gvi=gvi+1) begin: GEN_WWORD_LINE
    assign wword_line[gvi] = wr & (waddr == gvi[AW-1:0]);
  end 
  endgenerate
  generate
  for (gvi=0; gvi<DP; gvi=gvi+1) begin: GEN_MEN
  e603_subsys_gnrl_mem_line #(.DW(DW)) 
  U_mem_line (
  .clk(wclk), 
  .rst_n(wrst_n), 
  .wr(wword_line[gvi]), 
  .wdata(wdata), 
  .mem(mem[gvi*DW+DW-1:gvi*DW])
  );
  end 
  endgenerate
  e603_subsys_gnrl_data_mux #(.DW(DW), .N(DP))
  U_rdata_mux (
  .out_data(rdata_int),
  .in_data(mem),
  .sel(raddr)
  );
  generate
  if (REG_OUT > 0) begin: REG_OUT_1
e603_subsys_gnrl_dfflr #(DW) rdata_dfflr (rd, rdata_int, rdata, rclk, rrst_n);// VPP_NO_REG_PARSE
  end 
  else begin: REG_OUT_0
    assign rdata = rdata_int;
  end 
  endgenerate
endmodule 
module e603_subsys_gnrl_async_sdp_ram #(
  parameter DW = 8,
  parameter DP = 4,
  parameter DP_PTR_W = 2,
  parameter REG_OUT = 1,
  parameter PAYLOAD_NORST = 0,
  parameter AW = (DP <= 1) ? 1 : DP_PTR_W
)(
  input           wclk,
  input           wrst_n,
  input           wr,
  input  [AW-1:0] waddr,
  input  [DW-1:0] wdata,
  input           rclk,
  input           rrst_n,
  input           rd,
  input  [AW-1:0] raddr,
  output [DW-1:0] rdata
);
  wire    [DP-1:0] wword_line, rword_line;
  wire [DP*DW-1:0] mem;
  wire    [DW-1:0] rdata_int;
  genvar gvi;
  generate
  for (gvi=0; gvi<DP; gvi=gvi+1) begin: GEN_WWORD_LINE
    assign wword_line[gvi] = wr & (waddr == gvi[AW-1:0]);
  end 
  endgenerate
  generate
  for (gvi=0; gvi<DP; gvi=gvi+1) begin: GEN_MEN
  e603_subsys_gnrl_async_mem_line #(.DW(DW), .PAYLOAD_NORST(PAYLOAD_NORST)) 
  U_mem_line (
  .clk(wclk), 
  .rst_n(wrst_n), 
  .wr(wword_line[gvi]), 
  .wdata(wdata), 
  .mem(mem[gvi*DW+DW-1:gvi*DW])
  );
  end 
  endgenerate
  e603_subsys_gnrl_data_mux #(.DW(DW), .N(DP))
  U_rdata_mux (
  .out_data(rdata_int),
  .in_data(mem),
  .sel(raddr)
  );
  generate
  if (REG_OUT > 0) begin: REG_OUT_1
    if(PAYLOAD_NORST == 1) begin: payload_norst
    e603_subsys_gnrl_cdc_dffl  #(DW) rdata_gnrl_cdc_dest_dffl  (rd, rdata_int, rdata, rclk, rrst_n);// VPP_NO_REG_PARSE
    end
    else begin: payload_rst
    e603_subsys_gnrl_cdc_dfflr #(DW) rdata_gnrl_cdc_dest_dfflr (rd, rdata_int, rdata, rclk, rrst_n);// VPP_NO_REG_PARSE
    end
  end 
  else begin: REG_OUT_0
    assign rdata = rdata_int;
  end 
  endgenerate
endmodule 
`include "global.v"
module e603_subsys_gnrl_0dfflr # (
  parameter DW = 32
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
assign qout = dnxt;
endmodule
module e603_subsys_gnrl_0dffl # (
  parameter DW = 32
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk
);
assign qout = dnxt;
endmodule
module e603_subsys_gnrl_dfflrs # (
  parameter DW   = 32
, parameter [DW-1:0]  RST  = {DW{1'b1}}
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= RST;
  else if (lden == 1'b1)
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_cdc_dfflrs # (
  parameter DW   = 32
, parameter [DW-1:0]  RST  = {DW{1'b1}}
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= RST;
  else if (lden == 1'b1)
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_prot_dfflrs # (
  parameter DW   = 32
, parameter [DW-1:0]  RST  = {DW{1'b1}}
) (
  output              error,
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
localparam [0:0]    PAR_RESET   = (^RST) & 1;
reg [DW:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {PAR_RESET, RST};
  else if (lden == 1'b1)
    qout_r <= {^dnxt, dnxt};
end
assign qout = qout_r[DW-1:0];
assign error = qout_r[DW] != (^qout);
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_prot_cdc_dfflrs # (
  parameter DW   = 32
, parameter [DW-1:0]  RST  = {DW{1'b1}}
) (
  output              error,
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
localparam [0:0]    PAR_RESET   = (^RST) & 1;
reg [DW:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {PAR_RESET, RST};
  else if (lden == 1'b1)
    qout_r <= {^dnxt, dnxt};
end
assign qout = qout_r[DW-1:0];
assign error = qout_r[DW] != (^qout);
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_dfflr # (
  parameter DW   = 32
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else if (lden == 1'b1)
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_cdc_dfflr # (
  parameter DW   = 32
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else if (lden == 1'b1)
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_prot_dfflr # (
  parameter DW   = 32
) (
  output              error,
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {(DW+1){1'b0}};
  else if (lden == 1'b1)
    qout_r <= {^dnxt, dnxt};
end
assign qout = qout_r[DW-1:0];
assign error = qout_r[DW] != (^qout);
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_prot_cdc_dfflr # (
  parameter DW   = 32
) (
  output              error,
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {(DW+1){1'b0}};
  else if (lden == 1'b1)
    qout_r <= {^dnxt, dnxt};
end
assign qout = qout_r[DW-1:0];
assign error = qout_r[DW] != (^qout);
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_dfflrc # (
  parameter DW   = 32
) (
  input               clr,
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else if (clr == 1'b1)
    qout_r <= {DW{1'b0}};
  else if (lden == 1'b1)
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_cdc_dfflrc # (
  parameter DW   = 32
) (
  input               clr,
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else if (clr == 1'b1)
    qout_r <= {DW{1'b0}};
  else if (lden == 1'b1)
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_dffl # (
  parameter DW   = 32
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
// spyglass disable_block STARC-2.3.4.3
// SMD: Checks flip-flop asynchronous set or asynchronous reset
always @(posedge clk)
begin : DFF_PROC
  if (lden == 1'b1)
    qout_r <= dnxt;
end
// spyglass enable_block STARC-2.3.4.3
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_cdc_dffl # (
  parameter DW   = 32
) (
  input               lden,
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
// spyglass disable_block STARC-2.3.4.3
// SMD: Checks flip-flop asynchronous set or asynchronous reset
always @(posedge clk)
begin : DFF_PROC
  if (lden == 1'b1)
    qout_r <= dnxt;
end
// spyglass enable_block STARC-2.3.4.3
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_dff # (
  parameter DW   = 32
) (
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
// spyglass disable_block STARC-2.3.4.3
// SMD: Checks flip-flop asynchronous set or asynchronous reset
always @(posedge clk)
begin : DFF_PROC
    qout_r <= dnxt;
end
// spyglass enable_block STARC-2.3.4.3
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_cdc_dff # (
  parameter DW   = 32
) (
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
// spyglass disable_block STARC-2.3.4.3
// SMD: Checks flip-flop asynchronous set or asynchronous reset
always @(posedge clk)
begin : DFF_PROC
    qout_r <= dnxt;
end
// spyglass enable_block STARC-2.3.4.3
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_dffrs # (
  parameter DW   = 32
, parameter [DW-1:0]  RST  = {DW{1'b1}}
) (
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= RST;
  else
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_cdc_dffrs # (
  parameter DW   = 32
, parameter [DW-1:0]  RST  = {DW{1'b1}}
) (
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= RST;
  else
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
module e603_subsys_gnrl_dffr # (
  parameter DW   = 32
) (
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
endmodule
module e603_subsys_gnrl_cdc_dffr # (
  parameter DW   = 32
) (
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,
  input               clk,
  input               rst_n
);
reg [DW-1:0] qout_r;
// spyglass disable_block Ac_unsync01
// SMD: Checks unsynchronized crossings for scalar signals
// spyglass disable_block Ac_unsync02
// SMD: Checks unsynchronized crossings for vector signals
// spyglass disable_block Ar_asyncdeassert01
// SMD: Reports if reset signal is asynchronously deasserted
// spyglass disable_block Ar_unsync01
// SMD: Reports unsynchronized reset signals in the design
// spyglass disable_block Reset_sync02
// SMD: Reports asynchronous reset signals which are generated in asynchronous clock domain
// spyglass disable_block Ac_glitch04
// SMD: Reports clock domain crossings subject to glitches
// spyglass disable_block Clock_sync05a
// SMD: Reports primary inputs sampled by multiple clock domains
// spyglass disable_block Reset_sync04
// SMD: Reports asynchronous resets synchronized more than once in the same clock domain
// spyglass disable_block Ac_cdc01a
// SMD: Checks data loss for multi-flop or sync cell or qualifier synchronized clock domain
// SJ:  CDC register does not need to check for CDC rules
// spyglass disable_block UnrecSynthDir-ML 
// SMD: Synthesis directive is not recognized 
// SJ:  infer_multibit is okay to be here
always @(posedge clk or negedge rst_n)
begin : DFF_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else
    qout_r <= dnxt;
end
assign qout = qout_r[DW-1:0];
// spyglass enable_block UnrecSynthDir-ML
// spyglass enable_block Ac_unsync01
// spyglass enable_block Ac_unsync02
// spyglass enable_block Ar_asyncdeassert01
// spyglass enable_block Ar_unsync01
// spyglass enable_block Reset_sync02
// spyglass enable_block Ac_glitch04
// spyglass enable_block Clock_sync05a
// spyglass enable_block Reset_sync04
// spyglass enable_block Ac_cdc01a
endmodule
`include "global.v"
`include "global.v"
module e603_subsys_gnrl_fifo # (
  parameter CUT_READY = 0,
  parameter MSKO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter REGOUT_NORST = 0,
  parameter REG_OUT = 0,
  parameter DP   = 8,
  parameter DW   = 32
) (
  input           i_vld, 
  output          i_rdy, 
  input  [DW-1:0] i_dat,
  output          o_vld, 
  input           o_rdy, 
  output [DW-1:0] o_dat,
  input           clk,
  input           rst_n
);
genvar i;
generate 
  if(DP == 0) begin: gen_dp_eq1
     assign o_vld = i_vld;
     assign i_rdy = o_rdy;
     assign o_dat = i_dat;
  end
  else begin: gen_dp_gt0
    wire [DW-1:0] fifo_rf_din [DP-1:0];
    wire [DW-1:0] fifo_rf_r [DP-1:0];
    wire [DP-1:0] fifo_rf_en;
    wire wen = i_vld & i_rdy;
    wire ren = o_vld & o_rdy;
    wire [DP-1:0] rptr_vec_nxt; 
    wire [DP-1:0] rptr_vec_r;
    wire [DP-1:0] wptr_vec_nxt; 
    wire [DP-1:0] wptr_vec_r;
    if(DP == 1) begin:gen_rptr_dp_1
      assign rptr_vec_nxt = 1'b1; 
    end
    else begin:gen_rptr_dp_not_1
      assign rptr_vec_nxt = 
          rptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                          (rptr_vec_r << 1);
   end
    if(DP == 1) begin:gen_wptr_dp_1
      assign wptr_vec_nxt = 1'b1; 
    end
    else begin:gen_wptr_dp_not_1
      assign wptr_vec_nxt =
          wptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                          (wptr_vec_r << 1);
    end
// spyglass disable_block FlopSRConst
// SMD: master RTL_FDPE) is always set
// SJ:  Here is not a real issue
e603_subsys_gnrl_dfflrs #(1)    rptr_vec_0_dfflrs  (ren, rptr_vec_nxt[0]     , rptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflrs #(1)    wptr_vec_0_dfflrs  (wen, wptr_vec_nxt[0]     , wptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
// spyglass enable_block FlopSRConst
    if(DP > 1) begin:gen_dp_gt1
e603_subsys_gnrl_dfflr  #(DP-1) rptr_vec_31_dfflr  (ren, rptr_vec_nxt[DP-1:1], rptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP-1) wptr_vec_31_dfflr  (wen, wptr_vec_nxt[DP-1:1], wptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
    end
    wire [DP-1:0] i_vec;
    wire [DP-1:0] o_vec;
    wire [DP-1:0] vec_nxt; 
    wire [DP-1:0] vec_r;
    wire vec_en = (ren ^ wen );
e603_subsys_gnrl_dfflr  #(DP) vec_dfflr     (vec_en, vec_nxt, vec_r,     clk, rst_n);// VPP_NO_REG_PARSE
    assign i_vec = vec_r;
    assign o_vec = vec_r;
    if(DP == 1) begin:gen_cut_dp_eq1
        assign vec_nxt = wen ? 1'b1 : (vec_r >> 1);  
        if(CUT_READY == 1) begin:gen_cut_ready
          assign i_rdy = (~i_vec[DP-1]);
        end
        else begin:gen_no_cut_ready
          assign i_rdy = (~i_vec[DP-1]) | ren;
        end
    end
    else begin : no_cut_dp_gt1
      assign vec_nxt = wen ? {vec_r[DP-2:0], 1'b1} : (vec_r >> 1);  
      assign i_rdy = (~i_vec[DP-1]);
    end
    for (i=0; i<DP; i=i+1) begin:gen_fifo_rf
      assign fifo_rf_en[i] = wen & wptr_vec_r[i];
    if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_dffl  #(DW) fifo_rf_dffl (fifo_rf_en[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
    else begin: rst_gen
e603_subsys_gnrl_dfflr  #(DW) fifo_rf_dfflr (fifo_rf_en[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
      assign fifo_rf_din[i] = fifo_rf_en[i] ? i_dat : fifo_rf_r[i];
    end
    integer j;
    wire [DW-1:0] mux_rdat;
    if(REG_OUT == 0) begin:gen_rdat_output
    reg [DW-1:0] mux_rdat_t;
        always @*
        begin : rd_port_PROC
          mux_rdat_t = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_t = mux_rdat_t | ({DW{rptr_vec_r[j]}} & fifo_rf_r[j]);
          end
        end
    assign mux_rdat = mux_rdat_t;
    end
    else begin:gen_rdat_flp_output
        reg [DW-1:0] mux_rdat_rf_r;
        always @*
        begin : rd_port_PROC
          mux_rdat_rf_r = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_rf_r = mux_rdat_rf_r | ({DW{rptr_vec_nxt[j]}} & fifo_rf_r[j]);
          end
        end
        wire mux_rdat_ena = 
                        o_vld ? ren & vec_nxt[0] :
                                wen;
        wire [DW-1:0] mux_rdat_din = ~o_vec[1] ? i_dat : mux_rdat_rf_r;
      if(REGOUT_NORST == 0) begin:gen_rdat_output
e603_subsys_gnrl_dfflr #(DW) mux_rdat_dfflr  (mux_rdat_ena, mux_rdat_din, mux_rdat, clk, rst_n);// VPP_NO_REG_PARSE
      end
      else begin: gen_rdat_output_norst
e603_subsys_gnrl_dffl  #(DW) mux_rdat_dffl   (mux_rdat_ena, mux_rdat_din, mux_rdat, clk, rst_n);// VPP_NO_REG_PARSE
      end
`ifndef FPGA_SOURCE
`ifndef SYNTHESIS
        wire [DP-1:0] rptr_vec_din = ren ? rptr_vec_nxt : rptr_vec_r;
        wire [DW-1:0] mux_rdat_gold;
        reg [DW-1:0] mux_rdat_din_gold;
        always @*
        begin : rd_port_gold
          mux_rdat_din_gold = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_din_gold = mux_rdat_din_gold | ({DW{rptr_vec_din[j]}} & fifo_rf_din[j]);
          end
        end
e603_subsys_gnrl_dfflr #(DW) mux_rdat_gold_dfflr(mux_rdat_ena, mux_rdat_din_gold, mux_rdat_gold, clk, rst_n);// VPP_NO_REG_PARSE
`endif
`endif
    end
    if(MSKO == 1) begin:gen_mask_output
        assign o_dat = {DW{o_vld}} & mux_rdat;
    end
    else begin:gen_no_mask_output
        assign o_dat = mux_rdat;
    end
    assign o_vld = (o_vec[0]);
  end
endgenerate
endmodule 
module e603_subsys_gnrl_fifo_extends # (
  parameter CUT_READY = 0,
  parameter MSKO = 0,
  parameter PAYLOAD_NORST = 0,
  parameter REGOUT_NORST = 0,
  parameter REG_OUT = 0,
  parameter DP   = 8,
  parameter DW   = 32
) (
  input           i_vld, 
  output          i_rdy, 
  input  [DW-1:0] i_dat,
  output          o_vld, 
  input           o_rdy, 
  output [DW-1:0] o_dat,
  input           clk,
  input           rst_n
);
genvar i;
generate 
  if(DP == 0) begin: gen_dp_eq1
     assign o_vld = i_vld;
     assign i_rdy = o_rdy;
     assign o_dat = i_dat;
  end
  else begin: gen_dp_gt0
    wire [DW-1:0] fifo_rf_din [DP-1:0];
    wire [DW-1:0] fifo_rf_r [DP-1:0];
    wire [DP-1:0] fifo_rf_en;
    wire wen = i_vld & i_rdy;
    wire ren = o_vld & o_rdy;
    wire [DP-1:0] rptr_vec_din; 
    wire [DP-1:0] rptr_vec_nxt; 
    wire [DP-1:0] rptr_vec_r;
    wire [DP-1:0] wptr_vec_nxt; 
    wire [DP-1:0] wptr_vec_r;
    if(DP == 1) begin:gen_rptr_dp_1
      assign rptr_vec_nxt = 1'b1; 
    end
    else begin:gen_rptr_dp_not_1
      assign rptr_vec_nxt = 
          rptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                          (rptr_vec_r << 1);
   end
    if(DP == 1) begin:gen_wptr_dp_1
      assign wptr_vec_nxt = 1'b1; 
    end
    else begin:gen_wptr_dp_not_1
      assign wptr_vec_nxt =
          wptr_vec_r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                          (wptr_vec_r << 1);
    end
e603_subsys_gnrl_dfflrs #(1)    rptr_vec_0_dfflrs  (ren, rptr_vec_nxt[0]     , rptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflrs #(1)    wptr_vec_0_dfflrs  (wen, wptr_vec_nxt[0]     , wptr_vec_r[0]     , clk, rst_n);// VPP_NO_REG_PARSE
    if(DP > 1) begin:gen_dp_gt1
e603_subsys_gnrl_dfflr  #(DP-1) rptr_vec_31_dfflr  (ren, rptr_vec_nxt[DP-1:1], rptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
e603_subsys_gnrl_dfflr  #(DP-1) wptr_vec_31_dfflr  (wen, wptr_vec_nxt[DP-1:1], wptr_vec_r[DP-1:1], clk, rst_n);// VPP_NO_REG_PARSE
    end
    assign rptr_vec_din = ren ? rptr_vec_nxt : rptr_vec_r;
    wire [DP-1:0] i_vec;
    wire [DP-1:0] o_vec;
    wire [DP-1:0] vec_nxt; 
    wire [DP-1:0] vec_r;
    wire vec_en = (ren ^ wen );
e603_subsys_gnrl_dfflr  #(DP) vec_dfflr     (vec_en, vec_nxt, vec_r,     clk, rst_n);// VPP_NO_REG_PARSE
    assign i_vec = vec_r;
    assign o_vec = vec_r;
    if(DP == 1) begin:gen_cut_dp_eq1
        assign vec_nxt = wen ? 1'b1 : (vec_r >> 1);  
        if(CUT_READY == 1) begin:gen_cut_ready
          assign i_rdy = (~i_vec[DP-1]);
        end
        else begin:gen_no_cut_ready
          assign i_rdy = (~i_vec[DP-1]) | ren;
        end
    end
    else begin : no_cut_dp_gt1
      assign vec_nxt = wen ? {vec_r[DP-2:0], 1'b1} : (vec_r >> 1);  
     if(CUT_READY == 1) begin:gen_cut_ready_dp 
      assign i_rdy = (~i_vec[DP-1]);
     end
     else begin:gen_no_cut_ready_dp
      assign i_rdy = (~i_vec[DP-1]) | ren;
     end
    end
    for (i=0; i<DP; i=i+1) begin:gen_fifo_rf
      assign fifo_rf_en[i] = wen & wptr_vec_r[i];
    if(PAYLOAD_NORST == 1) begin:no_rst_gen
e603_subsys_gnrl_dffl  #(DW) fifo_rf_dffl (fifo_rf_en[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
    else begin: rst_gen
e603_subsys_gnrl_dfflr  #(DW) fifo_rf_dfflr (fifo_rf_en[i], i_dat, fifo_rf_r[i], clk, rst_n);// VPP_NO_REG_PARSE
    end
      assign fifo_rf_din[i] = fifo_rf_en[i] ? i_dat : fifo_rf_r[i];
    end
    integer j;
    wire [DW-1:0] mux_rdat;
    if(REG_OUT == 0) begin:gen_rdat_output
    reg [DW-1:0] mux_rdat_t;
        always @*
        begin : rd_port_PROC
          mux_rdat_t = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_t = mux_rdat_t | ({DW{rptr_vec_r[j]}} & fifo_rf_r[j]);
          end
        end
    assign mux_rdat = mux_rdat_t;
    end
    else begin:gen_rdat_flp_output
        reg [DW-1:0] mux_rdat_din;
        always @*
        begin : rd_port_PROC
          mux_rdat_din = {DW{1'b0}};
          for(j=0; j<DP; j=j+1) begin
            mux_rdat_din = mux_rdat_din | ({DW{rptr_vec_din[j]}} & fifo_rf_din[j]);
          end
        end
        wire mux_rdat_ena = 
                     (~o_vld) ? wen :
                     (vec_nxt[0] & ren);
e603_subsys_gnrl_dfflr #(DW) mux_rdat_dfflr  (mux_rdat_ena, mux_rdat_din, mux_rdat, clk, rst_n);// VPP_NO_REG_PARSE
    end
    if(MSKO == 1) begin:gen_mask_output
        assign o_dat = {DW{o_vld}} & mux_rdat;
    end
    else begin:gen_no_mask_output
        assign o_dat = mux_rdat;
    end
    assign o_vld = (o_vec[0]);
  end
endgenerate
endmodule 
`include "global.v"
`include "global.v"
