 /*                                                                      
  *  Copyright (c) 2018-2025 Nuclei System Technology, Inc.       
  *  All rights reserved.                                                
  */                                                                     
`include "global.v"
module e603_subsys_srams(
  input                            clk,
  input  rst_icache_ram,
  input                                 icache_tag0_cs,  
  input                                 icache_tag0_we,  
  input  [8-1:0]  icache_tag0_addr, 
  input  [22-1:0]  icache_tag0_wdata,          
  output [22-1:0]  icache_tag0_rdata,
  input                        clk_icache_tag0,
  input                                 icache_data0_cs,  
  input                                 icache_data0_we,  
  input  [11-1:0] icache_data0_addr, 
  input  [64-1:0] icache_data0_wdata,          
  output [64-1:0] icache_data0_rdata,
  input                        clk_icache_data0,
  input                                 icache_tag1_cs,  
  input                                 icache_tag1_we,  
  input  [8-1:0]  icache_tag1_addr, 
  input  [22-1:0]  icache_tag1_wdata,          
  output [22-1:0]  icache_tag1_rdata,
  input                        clk_icache_tag1,
  input                                 icache_data1_cs,  
  input                                 icache_data1_we,  
  input  [11-1:0] icache_data1_addr, 
  input  [64-1:0] icache_data1_wdata,          
  output [64-1:0] icache_data1_rdata,
  input                        clk_icache_data1,
  input  rst_dcache_ram,
  input                          clk_dcache_w0_tram,
  input                          clk_dcache_w1_tram,
  input                           dcache_w0_tram_cs,  
  input  [8-1:0]  dcache_w0_tram_addr,
  input                           dcache_w0_tram_we ,
  input  [21-1:0]  dcache_w0_tram_din,          
  output [21-1:0]  dcache_w0_tram_dout,
  input                           dcache_w1_tram_cs,  
  input  [8-1:0]  dcache_w1_tram_addr, 
  input                           dcache_w1_tram_we ,
  input  [21-1:0]  dcache_w1_tram_din,          
  output [21-1:0]  dcache_w1_tram_dout,
  input                          clk_dcache_dram_b0,
  input                           dcache_dram_b0_cs,  
  input                           dcache_dram_b0_we,  
  input  [10-1:0] dcache_dram_b0_addr, 
  input  [4-1:0] dcache_dram_b0_wem,
  input  [32-1:0] dcache_dram_b0_din,          
  output [32-1:0] dcache_dram_b0_dout,
  input                          clk_dcache_dram_b1,
  input                           dcache_dram_b1_cs,  
  input                           dcache_dram_b1_we,  
  input  [10-1:0] dcache_dram_b1_addr, 
  input  [4-1:0] dcache_dram_b1_wem,
  input  [32-1:0] dcache_dram_b1_din,          
  output [32-1:0] dcache_dram_b1_dout,
  input                          clk_dcache_dram_b2,
  input                           dcache_dram_b2_cs,  
  input                           dcache_dram_b2_we,  
  input  [10-1:0] dcache_dram_b2_addr, 
  input  [4-1:0] dcache_dram_b2_wem,
  input  [32-1:0] dcache_dram_b2_din,          
  output [32-1:0] dcache_dram_b2_dout,
  input                          clk_dcache_dram_b3,
  input                           dcache_dram_b3_cs,  
  input                           dcache_dram_b3_we,  
  input  [10-1:0] dcache_dram_b3_addr, 
  input  [4-1:0] dcache_dram_b3_wem,
  input  [32-1:0] dcache_dram_b3_din,          
  output [32-1:0] dcache_dram_b3_dout,
  input                          clk_dcache_dram_b4,
  input                           dcache_dram_b4_cs,  
  input                           dcache_dram_b4_we,  
  input  [10-1:0] dcache_dram_b4_addr, 
  input  [4-1:0] dcache_dram_b4_wem,
  input  [32-1:0] dcache_dram_b4_din,          
  output [32-1:0] dcache_dram_b4_dout,
  input                          clk_dcache_dram_b5,
  input                           dcache_dram_b5_cs,  
  input                           dcache_dram_b5_we,  
  input  [10-1:0] dcache_dram_b5_addr, 
  input  [4-1:0] dcache_dram_b5_wem,
  input  [32-1:0] dcache_dram_b5_din,          
  output [32-1:0] dcache_dram_b5_dout,
  input                          clk_dcache_dram_b6,
  input                           dcache_dram_b6_cs,  
  input                           dcache_dram_b6_we,  
  input  [10-1:0] dcache_dram_b6_addr, 
  input  [4-1:0] dcache_dram_b6_wem,
  input  [32-1:0] dcache_dram_b6_din,          
  output [32-1:0] dcache_dram_b6_dout,
  input                          clk_dcache_dram_b7,
  input                           dcache_dram_b7_cs,  
  input                           dcache_dram_b7_we,  
  input  [10-1:0] dcache_dram_b7_addr, 
  input  [4-1:0] dcache_dram_b7_wem,
  input  [32-1:0] dcache_dram_b7_din,          
  output [32-1:0] dcache_dram_b7_dout,
    input                                           rst_tlb_ram,
    input                                          clk_mmu_tlb_way0, 
    input                                          tlb_tram_way0_cs,
    input                                          tlb_dram_way0_cs,
    input                                          tlb_tram_way0_we,
    input                                          tlb_dram_way0_we,
    input [40-1:0]         tlb_tram_way0_wdata,
    input [27-1:0]         tlb_dram_way0_wdata,
    output  [40-1:0]       tlb_tram_way0_dout,
    output  [27-1:0]       tlb_dram_way0_dout,
    input [7-1:0]              tlb_tram_way0_addr,
    input [7-1:0]              tlb_dram_way0_addr,
    input                                          clk_mmu_tlb_way1, 
    input                                          tlb_tram_way1_cs,
    input                                          tlb_dram_way1_cs,
    input                                          tlb_tram_way1_we,
    input                                          tlb_dram_way1_we,
    input [40-1:0]         tlb_tram_way1_wdata,
    input [27-1:0]         tlb_dram_way1_wdata,
    output  [40-1:0]       tlb_tram_way1_dout,
    output  [27-1:0]       tlb_dram_way1_dout,
    input [7-1:0]              tlb_tram_way1_addr,
    input [7-1:0]              tlb_dram_way1_addr,
    input                                         rst_bht_ram,
  input                                                     bht_ram_bank0_cs, 
  input [9-2-1:0]  bht_ram_bank0_addr,
  input                                                     bht_ram_bank0_we,
  input [4*4-1:0]                          bht_ram_bank0_wem,
  input [4*4-1:0]                          bht_ram_bank0_din,
  output [4*4-1:0]                         bht_ram_bank0_dout,
  input clk_bht_ram_bank0,
  input                                                     bht_ram_bank1_cs, 
  input [9-2-1:0]  bht_ram_bank1_addr,
  input                                                     bht_ram_bank1_we,
  input [4*4-1:0]                          bht_ram_bank1_wem,
  input [4*4-1:0]                          bht_ram_bank1_din,
  output [4*4-1:0]                         bht_ram_bank1_dout,
  input clk_bht_ram_bank1,
  input                                                     bht_ram_bank2_cs, 
  input [9-2-1:0]  bht_ram_bank2_addr,
  input                                                     bht_ram_bank2_we,
  input [4*4-1:0]                          bht_ram_bank2_wem,
  input [4*4-1:0]                          bht_ram_bank2_din,
  output [4*4-1:0]                         bht_ram_bank2_dout,
  input clk_bht_ram_bank2,
  input                                                     bht_ram_bank3_cs, 
  input [9-2-1:0]  bht_ram_bank3_addr,
  input                                                     bht_ram_bank3_we,
  input [4*4-1:0]                          bht_ram_bank3_wem,
  input [4*4-1:0]                          bht_ram_bank3_din,
  output [4*4-1:0]                         bht_ram_bank3_dout,
  input clk_bht_ram_bank3,
    input                                         rst_btb_ram,
  input                                                 btb_ram_bank0_cs, 
  input [7-2-1:0] btb_ram_bank0_addr,
  input                                                 btb_ram_bank0_we,
  input [140-1:0]                          btb_ram_bank0_wem,
  input [140-1:0]                          btb_ram_bank0_din,
  output [140-1:0]                         btb_ram_bank0_dout,
  input clk_btb_ram_bank0,
  input                                                 btb_ram_bank1_cs, 
  input [7-2-1:0] btb_ram_bank1_addr,
  input                                                 btb_ram_bank1_we,
  input [140-1:0]                          btb_ram_bank1_wem,
  input [140-1:0]                          btb_ram_bank1_din,
  output [140-1:0]                         btb_ram_bank1_dout,
  input clk_btb_ram_bank1,
  input                                                 btb_ram_bank2_cs, 
  input [7-2-1:0] btb_ram_bank2_addr,
  input                                                 btb_ram_bank2_we,
  input [140-1:0]                          btb_ram_bank2_wem,
  input [140-1:0]                          btb_ram_bank2_din,
  output [140-1:0]                         btb_ram_bank2_dout,
  input clk_btb_ram_bank2,
  input                                                 btb_ram_bank3_cs, 
  input [7-2-1:0] btb_ram_bank3_addr,
  input                                                 btb_ram_bank3_we,
  input [140-1:0]                          btb_ram_bank3_wem,
  input [140-1:0]                          btb_ram_bank3_din,
  output [140-1:0]                         btb_ram_bank3_dout,
  input clk_btb_ram_bank3,
  input  dummy
);
    e603_data_ram u_data_b0_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b0_cs  ),  
                   .addr (dcache_dram_b0_addr), 
                   .we   (dcache_dram_b0_we),
                   .wem  (dcache_dram_b0_wem ),
                   .din  (dcache_dram_b0_din ),          
                   .dout (dcache_dram_b0_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b0)
                   );
    e603_data_ram u_data_b1_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b1_cs  ),  
                   .addr (dcache_dram_b1_addr), 
                   .we   (dcache_dram_b1_we),
                   .wem  (dcache_dram_b1_wem ),
                   .din  (dcache_dram_b1_din ),          
                   .dout (dcache_dram_b1_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b1)
                   );
    e603_data_ram u_data_b2_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b2_cs  ),  
                   .addr (dcache_dram_b2_addr), 
                   .we   (dcache_dram_b2_we),
                   .wem  (dcache_dram_b2_wem ),
                   .din  (dcache_dram_b2_din ),          
                   .dout (dcache_dram_b2_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b2)
                   );
    e603_data_ram u_data_b3_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b3_cs  ),  
                   .addr (dcache_dram_b3_addr), 
                   .we   (dcache_dram_b3_we),
                   .wem  (dcache_dram_b3_wem ),
                   .din  (dcache_dram_b3_din ),          
                   .dout (dcache_dram_b3_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b3)
                   );
    e603_data_ram u_data_b4_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b4_cs  ),  
                   .addr (dcache_dram_b4_addr), 
                   .we   (dcache_dram_b4_we),
                   .wem  (dcache_dram_b4_wem ),
                   .din  (dcache_dram_b4_din ),          
                   .dout (dcache_dram_b4_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b4)
                   );
    e603_data_ram u_data_b5_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b5_cs  ),  
                   .addr (dcache_dram_b5_addr), 
                   .we   (dcache_dram_b5_we),
                   .wem  (dcache_dram_b5_wem ),
                   .din  (dcache_dram_b5_din ),          
                   .dout (dcache_dram_b5_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b5)
                   );
    e603_data_ram u_data_b6_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b6_cs  ),  
                   .addr (dcache_dram_b6_addr), 
                   .we   (dcache_dram_b6_we),
                   .wem  (dcache_dram_b6_wem ),
                   .din  (dcache_dram_b6_din ),          
                   .dout (dcache_dram_b6_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b6)
                   );
    e603_data_ram u_data_b7_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_dram_b7_cs  ),  
                   .addr (dcache_dram_b7_addr), 
                   .we   (dcache_dram_b7_we),
                   .wem  (dcache_dram_b7_wem ),
                   .din  (dcache_dram_b7_din ),          
                   .dout (dcache_dram_b7_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_dram_b7)
                   );
    e603_dtag_ram u_dtag_w0_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_w0_tram_cs  ),  
                   .addr (dcache_w0_tram_addr), 
                   .we   (dcache_w0_tram_we),
                   .wem  ({3{dcache_w0_tram_we}}),
                   .din  (dcache_w0_tram_din ),          
                   .dout (dcache_w0_tram_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_w0_tram)
                   );
     e603_dtag_ram u_dtag_w1_ram(
                   .sd  (1'b0),
                   .ds  (1'b0),
                   .ls  (1'b0),
                   .cs   (dcache_w1_tram_cs  ),  
                   .addr (dcache_w1_tram_addr), 
                   .we   (dcache_w1_tram_we),
                   .wem  ({3{dcache_w1_tram_we}}),
                   .din  (dcache_w1_tram_din ),          
                   .dout (dcache_w1_tram_dout),
                   .rst_n (rst_dcache_ram),
                   .clk (clk_dcache_w1_tram)
                   );
  e603_icache_tag_ram u_icache_w0_tram (
    .sd   (1'b0   ),
    .ds   (1'b0   ),
    .ls   (1'b0   ),
    .cs   (icache_tag0_cs   ),
    .addr (icache_tag0_addr ),
    .we   (icache_tag0_we   ),
    .wem  ({3{icache_tag0_we}}  ),
    .din  (icache_tag0_wdata  ),
    .dout (icache_tag0_rdata ),
    .rst_n(rst_icache_ram  ),
    .clk  (clk_icache_tag0  )
    );
  e603_icache_data_ram u_icache_w0_dram (
    .sd   (1'b0   ),
    .ds   (1'b0   ),
    .ls   (1'b0   ),
    .cs   (icache_data0_cs   ),
    .addr (icache_data0_addr ),
    .we   (icache_data0_we   ),
    .wem  ({8{icache_data0_we }} ),
    .din  (icache_data0_wdata  ),
    .dout (icache_data0_rdata ),
    .rst_n(rst_icache_ram  ),
    .clk  (clk_icache_data0  )
    );
  e603_icache_tag_ram u_icache_w1_tram (
    .sd   (1'b0   ),
    .ds   (1'b0   ),
    .ls   (1'b0   ),
    .cs   (icache_tag1_cs   ),
    .addr (icache_tag1_addr ),
    .we   (icache_tag1_we   ),
    .wem  ({3{icache_tag1_we}}  ),
    .din  (icache_tag1_wdata  ),
    .dout (icache_tag1_rdata ),
    .rst_n(rst_icache_ram  ),
    .clk  (clk_icache_tag1  )
    );
  e603_icache_data_ram u_icache_w1_dram (
    .sd   (1'b0   ),
    .ds   (1'b0   ),
    .ls   (1'b0   ),
    .cs   (icache_data1_cs   ),
    .addr (icache_data1_addr ),
    .we   (icache_data1_we   ),
    .wem  ({8{icache_data1_we }} ),
    .din  (icache_data1_wdata  ),
    .dout (icache_data1_rdata ),
    .rst_n(rst_icache_ram  ),
    .clk  (clk_icache_data1  )
    );
  e603_tlb_tag_ram  u_tlb_ram_way0_tag (
        .sd     (1'b0   ),
        .ds     (1'b0   ),
        .ls     (1'b0   ),
        .cs     (tlb_tram_way0_cs),
        .we     (tlb_tram_way0_we),
        .wem    ({5{tlb_tram_way0_we}}),
        .addr   (tlb_tram_way0_addr),
        .din    (tlb_tram_way0_wdata),
        .dout   (tlb_tram_way0_dout),
        .rst_n  (rst_tlb_ram),
        .clk    (clk_mmu_tlb_way0)
    );
      e603_tlb_data_ram  u_tlb_ram_way0_data (
        .sd     (1'b0   ),
        .ds     (1'b0   ),
        .ls     (1'b0   ),
        .cs     (tlb_dram_way0_cs),
        .we     (tlb_dram_way0_we),
        .wem    ({4{tlb_dram_way0_we}}),
        .addr   (tlb_dram_way0_addr),
        .din    (tlb_dram_way0_wdata),
        .dout   (tlb_dram_way0_dout),
        .rst_n  (rst_tlb_ram),
        .clk    (clk_mmu_tlb_way0)
    );
  e603_tlb_tag_ram  u_tlb_ram_way1_tag (
        .sd     (1'b0   ),
        .ds     (1'b0   ),
        .ls     (1'b0   ),
        .cs     (tlb_tram_way1_cs),
        .we     (tlb_tram_way1_we),
        .wem    ({5{tlb_tram_way1_we}}),
        .addr   (tlb_tram_way1_addr),
        .din    (tlb_tram_way1_wdata),
        .dout   (tlb_tram_way1_dout),
        .rst_n  (rst_tlb_ram),
        .clk    (clk_mmu_tlb_way1)
    );
      e603_tlb_data_ram  u_tlb_ram_way1_data (
        .sd     (1'b0   ),
        .ds     (1'b0   ),
        .ls     (1'b0   ),
        .cs     (tlb_dram_way1_cs),
        .we     (tlb_dram_way1_we),
        .wem    ({4{tlb_dram_way1_we}}),
        .addr   (tlb_dram_way1_addr),
        .din    (tlb_dram_way1_wdata),
        .dout   (tlb_dram_way1_dout),
        .rst_n  (rst_tlb_ram),
        .clk    (clk_mmu_tlb_way1)
    );
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (512/4),
    .AW (9-2),
    .DW (4*4),
    .MW (4*4) 
)u_bht_ram_bank0 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_bht_ram),
    .we    (bht_ram_bank0_we),
    .clk   (clk_bht_ram_bank0),
    .din   (bht_ram_bank0_din),
    .addr  (bht_ram_bank0_addr),
    .cs    (bht_ram_bank0_cs),
    .wem   (bht_ram_bank0_wem),
    .dout  (bht_ram_bank0_dout)
);
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (512/4),
    .AW (9-2),
    .DW (4*4),
    .MW (4*4) 
)u_bht_ram_bank1 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_bht_ram),
    .we    (bht_ram_bank1_we),
    .clk   (clk_bht_ram_bank1),
    .din   (bht_ram_bank1_din),
    .addr  (bht_ram_bank1_addr),
    .cs    (bht_ram_bank1_cs),
    .wem   (bht_ram_bank1_wem),
    .dout  (bht_ram_bank1_dout)
);
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (512/4),
    .AW (9-2),
    .DW (4*4),
    .MW (4*4) 
)u_bht_ram_bank2 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_bht_ram),
    .we    (bht_ram_bank2_we),
    .clk   (clk_bht_ram_bank2),
    .din   (bht_ram_bank2_din),
    .addr  (bht_ram_bank2_addr),
    .cs    (bht_ram_bank2_cs),
    .wem   (bht_ram_bank2_wem),
    .dout  (bht_ram_bank2_dout)
);
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (512/4),
    .AW (9-2),
    .DW (4*4),
    .MW (4*4) 
)u_bht_ram_bank3 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_bht_ram),
    .we    (bht_ram_bank3_we),
    .clk   (clk_bht_ram_bank3),
    .din   (bht_ram_bank3_din),
    .addr  (bht_ram_bank3_addr),
    .cs    (bht_ram_bank3_cs),
    .wem   (bht_ram_bank3_wem),
    .dout  (bht_ram_bank3_dout)
);
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (32),
    .AW (7-2),
    .DW (140), 
    .MW (140) 
)u_btb_ram_bank0 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_btb_ram),
    .we    (btb_ram_bank0_we),
    .clk   (clk_btb_ram_bank0),
    .din   (btb_ram_bank0_din),
    .addr  (btb_ram_bank0_addr),
    .cs    (btb_ram_bank0_cs),
    .wem   (btb_ram_bank0_wem),
    .dout  (btb_ram_bank0_dout)
);
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (32),
    .AW (7-2),
    .DW (140), 
    .MW (140) 
)u_btb_ram_bank1 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_btb_ram),
    .we    (btb_ram_bank1_we),
    .clk   (clk_btb_ram_bank1),
    .din   (btb_ram_bank1_din),
    .addr  (btb_ram_bank1_addr),
    .cs    (btb_ram_bank1_cs),
    .wem   (btb_ram_bank1_wem),
    .dout  (btb_ram_bank1_dout)
);
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (32),
    .AW (7-2),
    .DW (140), 
    .MW (140) 
)u_btb_ram_bank2 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_btb_ram),
    .we    (btb_ram_bank2_we),
    .clk   (clk_btb_ram_bank2),
    .din   (btb_ram_bank2_din),
    .addr  (btb_ram_bank2_addr),
    .cs    (btb_ram_bank2_cs),
    .wem   (btb_ram_bank2_wem),
    .dout  (btb_ram_bank2_dout)
);
e603_gnrl_ram #(
    .FORCE_X2ZERO (1'b0),
    .DP (32),
    .AW (7-2),
    .DW (140), 
    .MW (140) 
)u_btb_ram_bank3 (
    .clkgate_bypass(1'b0),
    .sd    (1'b0),
    .ds    (1'b0),
    .ls    (1'b0),
    .rst_n (rst_btb_ram),
    .we    (btb_ram_bank3_we),
    .clk   (clk_btb_ram_bank3),
    .din   (btb_ram_bank3_din),
    .addr  (btb_ram_bank3_addr),
    .cs    (btb_ram_bank3_cs),
    .wem   (btb_ram_bank3_wem),
    .dout  (btb_ram_bank3_dout)
);
endmodule
