 /*                                                                      
  *  Copyright (c) 2018-2025 Nuclei System Technology, Inc.       
  *  All rights reserved.                                                
  */                                                                     
`include "global.v"
module soc_top #(
  parameter DDR_BG_WIDTH=1
)
(
  `ifdef DDR3_CONTROLLER
  inout  [31:0] ddr3_dq,
  inout  [3:0]  ddr3_dqs_n,
  inout  [3:0]  ddr3_dqs_p,
  output [13:0] ddr3_addr,
  output [2:0]  ddr3_ba,
  output        ddr3_ras_n,
  output        ddr3_cas_n,
  output        ddr3_we_n,
  output        ddr3_reset_n,
  output [0:0]  ddr3_ck_p,
  output [0:0]  ddr3_ck_n,
  output [0:0]  ddr3_cke,
  output [0:0]  ddr3_cs_n,
  output [3:0]  ddr3_dm,
  output [0:0]  ddr3_odt,
  output        init_calib_complete,
  input         ddr3_sys_clk_i,
  input         ddr3_sys_rst_i,
  `endif
  `ifdef DDR4_CONTROLLER
  inout  [7:0]  c0_ddr4_dm_dbi_n,
  inout  [63:0] c0_ddr4_dq,
  inout  [7:0]  c0_ddr4_dqs_c,
  inout  [7:0]  c0_ddr4_dqs_t,
  output        c0_ddr4_act_n,
  output [16:0] c0_ddr4_adr,
  output [1:0]  c0_ddr4_ba,
  output [DDR_BG_WIDTH-1:0]  c0_ddr4_bg,
  output [0:0]  c0_ddr4_cke,
  output [0:0]  c0_ddr4_odt,
  output [0:0]  c0_ddr4_cs_n,
  output [0:0]  c0_ddr4_ck_t,
  output [0:0]  c0_ddr4_ck_c,
  output        c0_ddr4_reset_n,
  output        init_calib_complete,
  input         ddr4_sys_clk_i,
  input         ddr4_sys_rst_i,
  `endif
  input              xec_sys_clk                   ,
  input              xmii_txc_i_ival               ,
  output             xmii_txc_o_oval               ,
  output             xmii_txc_o_oe                 ,
  input              gmii_rxc_i_ival               ,
  input              gmii_rxd_bit0_i_ival          ,
  output             gmii_txd_bit0_o_oval          ,
  input              gmii_rxd_bit1_i_ival          ,
  output             gmii_txd_bit1_o_oval          ,
  input              gmii_rxd_bit2_i_ival          ,
  output             gmii_txd_bit2_o_oval          ,
  input              gmii_rxd_bit3_i_ival          ,
  output             gmii_txd_bit3_o_oval          ,
  input              gmii_crs_i_ival               ,
  input              gmii_col_i_ival               ,
  input              gmii_rxdv_i_ival              ,
  input              gmii_rxer_i_ival              ,
  output             gmii_txen_o_oval              ,
  output             gmii_txer_o_oval              ,
  input              mdio_i_ival                   ,
  output             mdio_o_oval                   ,
  output             mdio_o_oe                     ,
  output             mdc_o_oval                    ,
  input   nex_clk,
  input   nex_rst_n,
  output  nex_o_clk,
  output [3:0] nex_o_data,
  input  por_rst_n,
  input  sys_rst_n,
  input  sys_clk,
`ifndef FPGA_SOURCE
  input  sys_clk_fast,
`endif
  input  aon_clk,
  input  evt_i,
  input  nmi_i,
  output core_wfi_mode,
  output core_sleep_value,
  input stop_on_reset,
  input   io_pads_jtag_TCK_i_ival,
  input   io_pads_jtag_TMS_i_ival,
  input   io_pads_jtag_TDI_i_ival,
  output  io_pads_jtag_TDO_o_oval,
  output  io_pads_jtag_tdo_drv_o_oval,
  output  io_pads_jtag_TMS_out_o_oval,
  output  io_pads_jtag_DRV_TMS_o_oval,
  output  io_pads_jtag_bk_o_oval     ,
  output  io_pads_qspi0_sck_o_oval,
  input   io_pads_qspi0_dq_0_i_ival,
  output  io_pads_qspi0_dq_0_o_oval,
  output  io_pads_qspi0_dq_0_o_oe,
  output  io_pads_qspi0_dq_0_o_ie,
  output  io_pads_qspi0_dq_0_o_pue,
  output  io_pads_qspi0_dq_0_o_ds,
  input   io_pads_qspi0_dq_1_i_ival,
  output  io_pads_qspi0_dq_1_o_oval,
  output  io_pads_qspi0_dq_1_o_oe,
  output  io_pads_qspi0_dq_1_o_ie,
  output  io_pads_qspi0_dq_1_o_pue,
  output  io_pads_qspi0_dq_1_o_ds,
  input   io_pads_qspi0_dq_2_i_ival,
  output  io_pads_qspi0_dq_2_o_oval,
  output  io_pads_qspi0_dq_2_o_oe,
  output  io_pads_qspi0_dq_2_o_ie,
  output  io_pads_qspi0_dq_2_o_pue,
  output  io_pads_qspi0_dq_2_o_ds,
  input   io_pads_qspi0_dq_3_i_ival,
  output  io_pads_qspi0_dq_3_o_oval,
  output  io_pads_qspi0_dq_3_o_oe,
  output  io_pads_qspi0_dq_3_o_ie,
  output  io_pads_qspi0_dq_3_o_pue,
  output  io_pads_qspi0_dq_3_o_ds,
  output  io_pads_qspi0_cs_0_o_oval,
  output  io_pads_qspi1_sck_o_oval,
  input   io_pads_qspi1_dq_0_i_ival,
  output  io_pads_qspi1_dq_0_o_oval,
  output  io_pads_qspi1_dq_0_o_oe,
  output  io_pads_qspi1_dq_0_o_ie,
  output  io_pads_qspi1_dq_0_o_pue,
  output  io_pads_qspi1_dq_0_o_ds,
  input   io_pads_qspi1_dq_1_i_ival,
  output  io_pads_qspi1_dq_1_o_oval,
  output  io_pads_qspi1_dq_1_o_oe,
  output  io_pads_qspi1_dq_1_o_ie,
  output  io_pads_qspi1_dq_1_o_pue,
  output  io_pads_qspi1_dq_1_o_ds,
  input   io_pads_qspi1_dq_2_i_ival,
  output  io_pads_qspi1_dq_2_o_oval,
  output  io_pads_qspi1_dq_2_o_oe,
  output  io_pads_qspi1_dq_2_o_ie,
  output  io_pads_qspi1_dq_2_o_pue,
  output  io_pads_qspi1_dq_2_o_ds,
  input   io_pads_qspi1_dq_3_i_ival,
  output  io_pads_qspi1_dq_3_o_oval,
  output  io_pads_qspi1_dq_3_o_oe,
  output  io_pads_qspi1_dq_3_o_ie,
  output  io_pads_qspi1_dq_3_o_pue,
  output  io_pads_qspi1_dq_3_o_ds,
  output  io_pads_qspi1_cs_0_o_oval,
  output  io_pads_qspi1_cs_1_o_oval,
  output  io_pads_qspi1_cs_2_o_oval,
  output  io_pads_qspi1_cs_3_o_oval,
  output  io_pads_qspi2_sck_o_oval,
  input   io_pads_qspi2_dq_0_i_ival,
  output  io_pads_qspi2_dq_0_o_oval,
  output  io_pads_qspi2_dq_0_o_oe,
  output  io_pads_qspi2_dq_0_o_ie,
  output  io_pads_qspi2_dq_0_o_pue,
  output  io_pads_qspi2_dq_0_o_ds,
  input   io_pads_qspi2_dq_1_i_ival,
  output  io_pads_qspi2_dq_1_o_oval,
  output  io_pads_qspi2_dq_1_o_oe,
  output  io_pads_qspi2_dq_1_o_ie,
  output  io_pads_qspi2_dq_1_o_pue,
  output  io_pads_qspi2_dq_1_o_ds,
  input   io_pads_qspi2_dq_2_i_ival,
  output  io_pads_qspi2_dq_2_o_oval,
  output  io_pads_qspi2_dq_2_o_oe,
  output  io_pads_qspi2_dq_2_o_ie,
  output  io_pads_qspi2_dq_2_o_pue,
  output  io_pads_qspi2_dq_2_o_ds,
  input   io_pads_qspi2_dq_3_i_ival,
  output  io_pads_qspi2_dq_3_o_oval,
  output  io_pads_qspi2_dq_3_o_oe,
  output  io_pads_qspi2_dq_3_o_ie,
  output  io_pads_qspi2_dq_3_o_pue,
  output  io_pads_qspi2_dq_3_o_ds,
  input   io_pads_qspi2_cs_0_i_ival,
  output  io_pads_qspi2_cs_0_o_oval,
  output  io_pads_qspi2_cs_0_o_oe,
  output  io_pads_qspi2_cs_0_o_ie,
  output  io_pads_qspi2_cs_0_o_pue,
  output  io_pads_qspi2_cs_0_o_ds,
  input   io_pads_uart0_rxd_i_ival,
  output  io_pads_uart0_rxd_o_oval,
  output  io_pads_uart0_rxd_o_oe,
  output  io_pads_uart0_rxd_o_ie,
  output  io_pads_uart0_rxd_o_pue,
  output  io_pads_uart0_rxd_o_ds,
  input   io_pads_uart0_txd_i_ival,
  output  io_pads_uart0_txd_o_oval,
  output  io_pads_uart0_txd_o_oe,
  output  io_pads_uart0_txd_o_ie,
  output  io_pads_uart0_txd_o_pue,
  output  io_pads_uart0_txd_o_ds
 );
 e603_subsys_top #(
    .DDR_BG_WIDTH(DDR_BG_WIDTH)
  ) 
  u_subsys_top(
  .por_rst_n(por_rst_n),
  .sys_rst_n(sys_rst_n),
  .sys_clk  (sys_clk  ),
`ifndef FPGA_SOURCE
  .sys_clk_fast(sys_clk_fast),
`endif
  .aon_clk  (aon_clk  ),
  .jtag_tdi                        (io_pads_jtag_TDI_i_ival),     
  .jtag_tdo                        (io_pads_jtag_TDO_o_oval),
  .jtag_tms                        (io_pads_jtag_TMS_i_ival),
  .jtag_tck                        (io_pads_jtag_TCK_i_ival),
  .jtag_tdo_drv                    (io_pads_jtag_tdo_drv_o_oval),
  .jtag_TMS_out                    (io_pads_jtag_TMS_out_o_oval),
  .jtag_DRV_TMS                    (io_pads_jtag_DRV_TMS_o_oval),
  .jtag_BK_TMS                     (io_pads_jtag_bk_o_oval     ),
   .nex_clk  (nex_clk),
   .nex_rst_n(nex_rst_n),
   .nex_o_clk(nex_o_clk),
   .nex_o_data  (nex_o_data),
  .test_mode(1'b0),
  .xec_sys_clk                   (xec_sys_clk                   ),
  .xmii_txc_i_ival               (xmii_txc_i_ival               ),
  .xmii_txc_o_oval               (xmii_txc_o_oval               ),
  .xmii_txc_o_oe                 (xmii_txc_o_oe                 ),
  .gmii_rxc_i_ival               (gmii_rxc_i_ival               ),
  .gmii_rxd_bit0_i_ival          (gmii_rxd_bit0_i_ival          ),
  .gmii_txd_bit0_o_oval          (gmii_txd_bit0_o_oval          ),
  .gmii_rxd_bit1_i_ival          (gmii_rxd_bit1_i_ival          ),
  .gmii_txd_bit1_o_oval          (gmii_txd_bit1_o_oval          ),
  .gmii_rxd_bit2_i_ival          (gmii_rxd_bit2_i_ival          ),
  .gmii_txd_bit2_o_oval          (gmii_txd_bit2_o_oval          ),
  .gmii_rxd_bit3_i_ival          (gmii_rxd_bit3_i_ival          ),
  .gmii_txd_bit3_o_oval          (gmii_txd_bit3_o_oval          ),
  .gmii_crs_i_ival               (gmii_crs_i_ival               ),
  .gmii_col_i_ival               (gmii_col_i_ival               ),
  .gmii_rxdv_i_ival              (gmii_rxdv_i_ival              ),
  .gmii_rxer_i_ival              (gmii_rxer_i_ival              ),
  .gmii_txen_o_oval              (gmii_txen_o_oval              ),
  .gmii_txer_o_oval              (gmii_txer_o_oval              ),
  .mdio_i_ival                   (mdio_i_ival                   ),
  .mdio_o_oval                   (mdio_o_oval                   ),
  .mdio_o_oe                     (mdio_o_oe                     ),
  .mdc_o_oval                    (mdc_o_oval                    ),
    .io_pads_qspi0_sck_i_ival (1'b1    ),
    .io_pads_qspi0_sck_o_oval (io_pads_qspi0_sck_o_oval    ),
    .io_pads_qspi0_sck_o_oe   (      ),
    .io_pads_qspi0_sck_o_ie   (      ),
    .io_pads_qspi0_sck_o_pue  (     ),
    .io_pads_qspi0_sck_o_ds   (      ),
    .io_pads_qspi0_dq_0_i_ival(io_pads_qspi0_dq_0_i_ival  & io_pads_qspi0_dq_0_o_ie ),
    .io_pads_qspi0_dq_0_o_oval(io_pads_qspi0_dq_0_o_oval   ),
    .io_pads_qspi0_dq_0_o_oe  (io_pads_qspi0_dq_0_o_oe     ),
    .io_pads_qspi0_dq_0_o_ie  (io_pads_qspi0_dq_0_o_ie     ),
    .io_pads_qspi0_dq_0_o_pue (io_pads_qspi0_dq_0_o_pue    ),
    .io_pads_qspi0_dq_0_o_ds  (io_pads_qspi0_dq_0_o_ds     ),
    .io_pads_qspi0_dq_1_i_ival(io_pads_qspi0_dq_1_i_ival & io_pads_qspi0_dq_1_o_ie ),
    .io_pads_qspi0_dq_1_o_oval(io_pads_qspi0_dq_1_o_oval   ),
    .io_pads_qspi0_dq_1_o_oe  (io_pads_qspi0_dq_1_o_oe     ),
    .io_pads_qspi0_dq_1_o_ie  (io_pads_qspi0_dq_1_o_ie     ),
    .io_pads_qspi0_dq_1_o_pue (io_pads_qspi0_dq_1_o_pue    ),
    .io_pads_qspi0_dq_1_o_ds  (io_pads_qspi0_dq_1_o_ds     ),
    .io_pads_qspi0_dq_2_i_ival(io_pads_qspi0_dq_2_i_ival & io_pads_qspi0_dq_2_o_ie  ),
    .io_pads_qspi0_dq_2_o_oval(io_pads_qspi0_dq_2_o_oval   ),
    .io_pads_qspi0_dq_2_o_oe  (io_pads_qspi0_dq_2_o_oe     ),
    .io_pads_qspi0_dq_2_o_ie  (io_pads_qspi0_dq_2_o_ie     ),
    .io_pads_qspi0_dq_2_o_pue (io_pads_qspi0_dq_2_o_pue    ),
    .io_pads_qspi0_dq_2_o_ds  (io_pads_qspi0_dq_2_o_ds     ),
    .io_pads_qspi0_dq_3_i_ival(io_pads_qspi0_dq_3_i_ival & io_pads_qspi0_dq_3_o_ie   ),
    .io_pads_qspi0_dq_3_o_oval(io_pads_qspi0_dq_3_o_oval   ),
    .io_pads_qspi0_dq_3_o_oe  (io_pads_qspi0_dq_3_o_oe     ),
    .io_pads_qspi0_dq_3_o_ie  (io_pads_qspi0_dq_3_o_ie     ),
    .io_pads_qspi0_dq_3_o_pue (io_pads_qspi0_dq_3_o_pue    ),
    .io_pads_qspi0_dq_3_o_ds  (io_pads_qspi0_dq_3_o_ds     ),
    .io_pads_qspi0_cs_0_i_ival(1'b1   ),
    .io_pads_qspi0_cs_0_o_oval(io_pads_qspi0_cs_0_o_oval   ),
    .io_pads_qspi0_cs_0_o_oe  (     ),
    .io_pads_qspi0_cs_0_o_ie  (     ),
    .io_pads_qspi0_cs_0_o_pue (    ),
    .io_pads_qspi0_cs_0_o_ds  (     ),
    .io_pads_qspi1_sck_i_ival (1'b1    ),
    .io_pads_qspi1_sck_o_oval (io_pads_qspi1_sck_o_oval    ),
    .io_pads_qspi1_sck_o_oe   (      ),
    .io_pads_qspi1_sck_o_ie   (      ),
    .io_pads_qspi1_sck_o_pue  (     ),
    .io_pads_qspi1_sck_o_ds   (      ),
    .io_pads_qspi1_dq_0_i_ival(io_pads_qspi1_dq_0_i_ival  & io_pads_qspi1_dq_0_o_ie ),
    .io_pads_qspi1_dq_0_o_oval(io_pads_qspi1_dq_0_o_oval   ),
    .io_pads_qspi1_dq_0_o_oe  (io_pads_qspi1_dq_0_o_oe     ),
    .io_pads_qspi1_dq_0_o_ie  (io_pads_qspi1_dq_0_o_ie     ),
    .io_pads_qspi1_dq_0_o_pue (io_pads_qspi1_dq_0_o_pue    ),
    .io_pads_qspi1_dq_0_o_ds  (io_pads_qspi1_dq_0_o_ds     ),
    .io_pads_qspi1_dq_1_i_ival(io_pads_qspi1_dq_1_i_ival & io_pads_qspi1_dq_1_o_ie ),
    .io_pads_qspi1_dq_1_o_oval(io_pads_qspi1_dq_1_o_oval   ),
    .io_pads_qspi1_dq_1_o_oe  (io_pads_qspi1_dq_1_o_oe     ),
    .io_pads_qspi1_dq_1_o_ie  (io_pads_qspi1_dq_1_o_ie     ),
    .io_pads_qspi1_dq_1_o_pue (io_pads_qspi1_dq_1_o_pue    ),
    .io_pads_qspi1_dq_1_o_ds  (io_pads_qspi1_dq_1_o_ds     ),
    .io_pads_qspi1_dq_2_i_ival(io_pads_qspi1_dq_2_i_ival & io_pads_qspi1_dq_2_o_ie  ),
    .io_pads_qspi1_dq_2_o_oval(io_pads_qspi1_dq_2_o_oval   ),
    .io_pads_qspi1_dq_2_o_oe  (io_pads_qspi1_dq_2_o_oe     ),
    .io_pads_qspi1_dq_2_o_ie  (io_pads_qspi1_dq_2_o_ie     ),
    .io_pads_qspi1_dq_2_o_pue (io_pads_qspi1_dq_2_o_pue    ),
    .io_pads_qspi1_dq_2_o_ds  (io_pads_qspi1_dq_2_o_ds     ),
    .io_pads_qspi1_dq_3_i_ival(io_pads_qspi1_dq_3_i_ival & io_pads_qspi1_dq_3_o_ie   ),
    .io_pads_qspi1_dq_3_o_oval(io_pads_qspi1_dq_3_o_oval   ),
    .io_pads_qspi1_dq_3_o_oe  (io_pads_qspi1_dq_3_o_oe     ),
    .io_pads_qspi1_dq_3_o_ie  (io_pads_qspi1_dq_3_o_ie     ),
    .io_pads_qspi1_dq_3_o_pue (io_pads_qspi1_dq_3_o_pue    ),
    .io_pads_qspi1_dq_3_o_ds  (io_pads_qspi1_dq_3_o_ds     ),
    .io_pads_qspi1_cs_0_i_ival(1'b1   ),
    .io_pads_qspi1_cs_0_o_oval(io_pads_qspi1_cs_0_o_oval   ),
    .io_pads_qspi1_cs_0_o_oe  (     ),
    .io_pads_qspi1_cs_0_o_ie  (     ),
    .io_pads_qspi1_cs_0_o_pue (    ),
    .io_pads_qspi1_cs_0_o_ds  (     ),
    .io_pads_qspi1_cs_1_i_ival(1'b1   ),
    .io_pads_qspi1_cs_1_o_oval(io_pads_qspi1_cs_1_o_oval   ),
    .io_pads_qspi1_cs_1_o_oe  (     ),
    .io_pads_qspi1_cs_1_o_ie  (     ),
    .io_pads_qspi1_cs_1_o_pue (    ),
    .io_pads_qspi1_cs_1_o_ds  (     ),
    .io_pads_qspi1_cs_2_i_ival(1'b1   ),
    .io_pads_qspi1_cs_2_o_oval(io_pads_qspi1_cs_2_o_oval   ),
    .io_pads_qspi1_cs_2_o_oe  (     ),
    .io_pads_qspi1_cs_2_o_ie  (     ),
    .io_pads_qspi1_cs_2_o_pue (    ),
    .io_pads_qspi1_cs_2_o_ds  (     ),
    .io_pads_qspi1_cs_3_i_ival(1'b1   ),
    .io_pads_qspi1_cs_3_o_oval(io_pads_qspi1_cs_3_o_oval   ),
    .io_pads_qspi1_cs_3_o_oe  (     ),
    .io_pads_qspi1_cs_3_o_ie  (     ),
    .io_pads_qspi1_cs_3_o_pue (    ),
    .io_pads_qspi1_cs_3_o_ds  (     ),
    .io_pads_qspi2_sck_i_ival (1'b1    ),
    .io_pads_qspi2_sck_o_oval (io_pads_qspi2_sck_o_oval    ),
    .io_pads_qspi2_sck_o_oe   (      ),
    .io_pads_qspi2_sck_o_ie   (      ),
    .io_pads_qspi2_sck_o_pue  (     ),
    .io_pads_qspi2_sck_o_ds   (      ),
    .io_pads_qspi2_dq_0_i_ival(io_pads_qspi2_dq_0_i_ival  & io_pads_qspi2_dq_0_o_ie ),
    .io_pads_qspi2_dq_0_o_oval(io_pads_qspi2_dq_0_o_oval   ),
    .io_pads_qspi2_dq_0_o_oe  (io_pads_qspi2_dq_0_o_oe     ),
    .io_pads_qspi2_dq_0_o_ie  (io_pads_qspi2_dq_0_o_ie     ),
    .io_pads_qspi2_dq_0_o_pue (io_pads_qspi2_dq_0_o_pue    ),
    .io_pads_qspi2_dq_0_o_ds  (io_pads_qspi2_dq_0_o_ds     ),
    .io_pads_qspi2_dq_1_i_ival(io_pads_qspi2_dq_1_i_ival & io_pads_qspi2_dq_1_o_ie ),
    .io_pads_qspi2_dq_1_o_oval(io_pads_qspi2_dq_1_o_oval   ),
    .io_pads_qspi2_dq_1_o_oe  (io_pads_qspi2_dq_1_o_oe     ),
    .io_pads_qspi2_dq_1_o_ie  (io_pads_qspi2_dq_1_o_ie     ),
    .io_pads_qspi2_dq_1_o_pue (io_pads_qspi2_dq_1_o_pue    ),
    .io_pads_qspi2_dq_1_o_ds  (io_pads_qspi2_dq_1_o_ds     ),
    .io_pads_qspi2_dq_2_i_ival(io_pads_qspi2_dq_2_i_ival & io_pads_qspi2_dq_2_o_ie  ),
    .io_pads_qspi2_dq_2_o_oval(io_pads_qspi2_dq_2_o_oval   ),
    .io_pads_qspi2_dq_2_o_oe  (io_pads_qspi2_dq_2_o_oe     ),
    .io_pads_qspi2_dq_2_o_ie  (io_pads_qspi2_dq_2_o_ie     ),
    .io_pads_qspi2_dq_2_o_pue (io_pads_qspi2_dq_2_o_pue    ),
    .io_pads_qspi2_dq_2_o_ds  (io_pads_qspi2_dq_2_o_ds     ),
    .io_pads_qspi2_dq_3_i_ival(io_pads_qspi2_dq_3_i_ival & io_pads_qspi2_dq_3_o_ie   ),
    .io_pads_qspi2_dq_3_o_oval(io_pads_qspi2_dq_3_o_oval   ),
    .io_pads_qspi2_dq_3_o_oe  (io_pads_qspi2_dq_3_o_oe     ),
    .io_pads_qspi2_dq_3_o_ie  (io_pads_qspi2_dq_3_o_ie     ),
    .io_pads_qspi2_dq_3_o_pue (io_pads_qspi2_dq_3_o_pue    ),
    .io_pads_qspi2_dq_3_o_ds  (io_pads_qspi2_dq_3_o_ds     ),
    .io_pads_qspi2_cs_0_i_ival(io_pads_qspi2_cs_0_i_ival   ),
    .io_pads_qspi2_cs_0_o_oval(io_pads_qspi2_cs_0_o_oval   ),
    .io_pads_qspi2_cs_0_o_oe  (io_pads_qspi2_cs_0_o_oe     ),
    .io_pads_qspi2_cs_0_o_ie  (io_pads_qspi2_cs_0_o_ie     ),
    .io_pads_qspi2_cs_0_o_pue (io_pads_qspi2_cs_0_o_pue    ),
    .io_pads_qspi2_cs_0_o_ds  (io_pads_qspi2_cs_0_o_ds     ),
    .io_pads_uart0_rxd_i_ival (io_pads_uart0_rxd_i_ival & io_pads_uart0_rxd_o_ie),
    .io_pads_uart0_rxd_o_oval (io_pads_uart0_rxd_o_oval),
    .io_pads_uart0_rxd_o_oe   (io_pads_uart0_rxd_o_oe),
    .io_pads_uart0_rxd_o_ie   (io_pads_uart0_rxd_o_ie),
    .io_pads_uart0_rxd_o_pue  (io_pads_uart0_rxd_o_pue),
    .io_pads_uart0_rxd_o_ds   (io_pads_uart0_rxd_o_ds),
    .io_pads_uart0_txd_i_ival (io_pads_uart0_txd_i_ival & io_pads_uart0_txd_o_ie),
    .io_pads_uart0_txd_o_oval (io_pads_uart0_txd_o_oval),
    .io_pads_uart0_txd_o_oe   (io_pads_uart0_txd_o_oe),
    .io_pads_uart0_txd_o_ie   (io_pads_uart0_txd_o_ie),
    .io_pads_uart0_txd_o_pue  (io_pads_uart0_txd_o_pue),
    .io_pads_uart0_txd_o_ds   (io_pads_uart0_txd_o_ds),
  `ifdef DDR3_CONTROLLER
  .ddr3_addr           (ddr3_addr),
  .ddr3_ba             (ddr3_ba),
  .ddr3_cas_n          (ddr3_cas_n),
  .ddr3_ck_n           (ddr3_ck_n),
  .ddr3_ck_p           (ddr3_ck_p),
  .ddr3_cke            (ddr3_cke),
  .ddr3_ras_n          (ddr3_ras_n),
  .ddr3_we_n           (ddr3_we_n),
  .ddr3_dq             (ddr3_dq),
  .ddr3_dqs_n          (ddr3_dqs_n),
  .ddr3_dqs_p          (ddr3_dqs_p),
  .ddr3_reset_n        (ddr3_reset_n),
  .ddr3_sys_clk_i      (ddr3_sys_clk_i),
  .ddr3_sys_rst_i      (ddr3_sys_rst_i),
  .ddr3_cs_n           (ddr3_cs_n),
  .ddr3_dm             (ddr3_dm),
  .ddr3_odt            (ddr3_odt),
  .init_calib_complete (init_calib_complete),
  `endif
  `ifdef DDR4_CONTROLLER
  .c0_ddr4_dm_dbi_n    (c0_ddr4_dm_dbi_n   ),
  .c0_ddr4_dq          (c0_ddr4_dq         ),
  .c0_ddr4_dqs_c       (c0_ddr4_dqs_c      ),
  .c0_ddr4_dqs_t       (c0_ddr4_dqs_t      ),
  .c0_ddr4_act_n       (c0_ddr4_act_n      ),
  .c0_ddr4_adr         (c0_ddr4_adr        ),
  .c0_ddr4_ba          (c0_ddr4_ba         ),
  .c0_ddr4_bg          (c0_ddr4_bg         ),
  .c0_ddr4_cke         (c0_ddr4_cke        ),
  .c0_ddr4_odt         (c0_ddr4_odt        ),
  .c0_ddr4_cs_n        (c0_ddr4_cs_n       ),
  .c0_ddr4_ck_t        (c0_ddr4_ck_t       ),
  .c0_ddr4_ck_c        (c0_ddr4_ck_c       ),
  .c0_ddr4_reset_n     (c0_ddr4_reset_n    ),
  .init_calib_complete (init_calib_complete),
  .ddr4_sys_clk_i      (ddr4_sys_clk_i      ),
  .ddr4_sys_rst_i      (ddr4_sys_rst_i     ),
  `endif
  `ifdef TEMAC_CONTROLLER
  .temac_axi_aclk    (temac_axi_aclk   ), 
  .temac_axi_aresetn (temac_axi_aresetn),
  .phy_tx_clk        (phy_tx_clk ),
  .phy_rx_clk        (phy_rx_clk ),
  .phy_crs           (phy_crs    ),
  .phy_dv            (phy_dv     ),
  .phy_rx_data       (phy_rx_data),
  .phy_col           (phy_col    ),
  .phy_rx_er         (phy_rx_er  ),
  .phy_rst_n         (phy_rst_n  ),
  .phy_tx_en         (phy_tx_en  ),
  .phy_tx_data       (phy_tx_data),
  .io_pins_mdio_i_ival (io_pins_mdio_i_ival  & io_pins_mdio_o_ie),
  .io_pins_mdio_o_oval (io_pins_mdio_o_oval  ),
  .io_pins_mdio_o_oe   (io_pins_mdio_o_oe    ),
  .io_pins_mdio_o_ie   (io_pins_mdio_o_ie    ),
  .io_pins_mdio_o_pue  (io_pins_mdio_o_pue   ),
  .io_pins_mdio_o_ds   (io_pins_mdio_o_ds    ),
  .phy_mdc           (phy_mdc    ),
  `endif
  .stop_on_reset    (stop_on_reset),
  .evt_i               (evt_i),
  .nmi_i               (nmi_i),
  .core_sleep_value    (core_sleep_value),
  .core_wfi_mode       (core_wfi_mode) 
  );
endmodule
